magic
tech gf180mcuD
magscale 1 5
timestamp 1701345104
<< obsm1 >>
rect 672 855 279328 248166
<< metal2 >>
rect 5488 0 5544 400
rect 6384 0 6440 400
rect 7280 0 7336 400
rect 8176 0 8232 400
rect 9072 0 9128 400
rect 9968 0 10024 400
rect 10864 0 10920 400
rect 11760 0 11816 400
rect 12656 0 12712 400
rect 13552 0 13608 400
rect 14448 0 14504 400
rect 15344 0 15400 400
rect 16240 0 16296 400
rect 17136 0 17192 400
rect 18032 0 18088 400
rect 18928 0 18984 400
rect 19824 0 19880 400
rect 20720 0 20776 400
rect 21616 0 21672 400
rect 22512 0 22568 400
rect 23408 0 23464 400
rect 24304 0 24360 400
rect 25200 0 25256 400
rect 26096 0 26152 400
rect 26992 0 27048 400
rect 27888 0 27944 400
rect 28784 0 28840 400
rect 29680 0 29736 400
rect 30576 0 30632 400
rect 31472 0 31528 400
rect 32368 0 32424 400
rect 33264 0 33320 400
rect 34160 0 34216 400
rect 35056 0 35112 400
rect 35952 0 36008 400
rect 36848 0 36904 400
rect 37744 0 37800 400
rect 38640 0 38696 400
rect 39536 0 39592 400
rect 40432 0 40488 400
rect 41328 0 41384 400
rect 42224 0 42280 400
rect 43120 0 43176 400
rect 44016 0 44072 400
rect 44912 0 44968 400
rect 45808 0 45864 400
rect 46704 0 46760 400
rect 47600 0 47656 400
rect 48496 0 48552 400
rect 49392 0 49448 400
rect 50288 0 50344 400
rect 51184 0 51240 400
rect 52080 0 52136 400
rect 52976 0 53032 400
rect 53872 0 53928 400
rect 54768 0 54824 400
rect 55664 0 55720 400
rect 56560 0 56616 400
rect 57456 0 57512 400
rect 58352 0 58408 400
rect 59248 0 59304 400
rect 60144 0 60200 400
rect 61040 0 61096 400
rect 61936 0 61992 400
rect 62832 0 62888 400
rect 63728 0 63784 400
rect 64624 0 64680 400
rect 65520 0 65576 400
rect 66416 0 66472 400
rect 67312 0 67368 400
rect 68208 0 68264 400
rect 69104 0 69160 400
rect 70000 0 70056 400
rect 70896 0 70952 400
rect 71792 0 71848 400
rect 72688 0 72744 400
rect 73584 0 73640 400
rect 74480 0 74536 400
rect 75376 0 75432 400
rect 76272 0 76328 400
rect 77168 0 77224 400
rect 78064 0 78120 400
rect 78960 0 79016 400
rect 79856 0 79912 400
rect 80752 0 80808 400
rect 81648 0 81704 400
rect 82544 0 82600 400
rect 83440 0 83496 400
rect 84336 0 84392 400
rect 85232 0 85288 400
rect 86128 0 86184 400
rect 87024 0 87080 400
rect 87920 0 87976 400
rect 88816 0 88872 400
rect 89712 0 89768 400
rect 90608 0 90664 400
rect 91504 0 91560 400
rect 92400 0 92456 400
rect 93296 0 93352 400
rect 94192 0 94248 400
rect 95088 0 95144 400
rect 95984 0 96040 400
rect 96880 0 96936 400
rect 97776 0 97832 400
rect 98672 0 98728 400
rect 99568 0 99624 400
rect 100464 0 100520 400
rect 101360 0 101416 400
rect 102256 0 102312 400
rect 103152 0 103208 400
rect 104048 0 104104 400
rect 104944 0 105000 400
rect 105840 0 105896 400
rect 106736 0 106792 400
rect 107632 0 107688 400
rect 108528 0 108584 400
rect 109424 0 109480 400
rect 110320 0 110376 400
rect 111216 0 111272 400
rect 112112 0 112168 400
rect 113008 0 113064 400
rect 113904 0 113960 400
rect 114800 0 114856 400
rect 115696 0 115752 400
rect 116592 0 116648 400
rect 117488 0 117544 400
rect 118384 0 118440 400
rect 119280 0 119336 400
rect 120176 0 120232 400
rect 121072 0 121128 400
rect 121968 0 122024 400
rect 122864 0 122920 400
rect 123760 0 123816 400
rect 124656 0 124712 400
rect 125552 0 125608 400
rect 126448 0 126504 400
rect 127344 0 127400 400
rect 128240 0 128296 400
rect 129136 0 129192 400
rect 130032 0 130088 400
rect 130928 0 130984 400
rect 131824 0 131880 400
rect 132720 0 132776 400
rect 133616 0 133672 400
rect 134512 0 134568 400
rect 135408 0 135464 400
rect 136304 0 136360 400
rect 137200 0 137256 400
rect 138096 0 138152 400
rect 138992 0 139048 400
rect 139888 0 139944 400
rect 140784 0 140840 400
rect 141680 0 141736 400
rect 142576 0 142632 400
rect 143472 0 143528 400
rect 144368 0 144424 400
rect 145264 0 145320 400
rect 146160 0 146216 400
rect 147056 0 147112 400
rect 147952 0 148008 400
rect 148848 0 148904 400
rect 149744 0 149800 400
rect 150640 0 150696 400
rect 151536 0 151592 400
rect 152432 0 152488 400
rect 153328 0 153384 400
rect 154224 0 154280 400
rect 155120 0 155176 400
rect 156016 0 156072 400
rect 156912 0 156968 400
rect 157808 0 157864 400
rect 158704 0 158760 400
rect 159600 0 159656 400
rect 160496 0 160552 400
rect 161392 0 161448 400
rect 162288 0 162344 400
rect 163184 0 163240 400
rect 164080 0 164136 400
rect 164976 0 165032 400
rect 165872 0 165928 400
rect 166768 0 166824 400
rect 167664 0 167720 400
rect 168560 0 168616 400
rect 169456 0 169512 400
rect 170352 0 170408 400
rect 171248 0 171304 400
rect 172144 0 172200 400
rect 173040 0 173096 400
rect 173936 0 173992 400
rect 174832 0 174888 400
rect 175728 0 175784 400
rect 176624 0 176680 400
rect 177520 0 177576 400
rect 178416 0 178472 400
rect 179312 0 179368 400
rect 180208 0 180264 400
rect 181104 0 181160 400
rect 182000 0 182056 400
rect 182896 0 182952 400
rect 183792 0 183848 400
rect 184688 0 184744 400
rect 185584 0 185640 400
rect 186480 0 186536 400
rect 187376 0 187432 400
rect 188272 0 188328 400
rect 189168 0 189224 400
rect 190064 0 190120 400
rect 190960 0 191016 400
rect 191856 0 191912 400
rect 192752 0 192808 400
rect 193648 0 193704 400
rect 194544 0 194600 400
rect 195440 0 195496 400
rect 196336 0 196392 400
rect 197232 0 197288 400
rect 198128 0 198184 400
rect 199024 0 199080 400
rect 199920 0 199976 400
rect 200816 0 200872 400
rect 201712 0 201768 400
rect 202608 0 202664 400
rect 203504 0 203560 400
rect 204400 0 204456 400
rect 205296 0 205352 400
rect 206192 0 206248 400
rect 207088 0 207144 400
rect 207984 0 208040 400
rect 208880 0 208936 400
rect 209776 0 209832 400
rect 210672 0 210728 400
rect 211568 0 211624 400
rect 212464 0 212520 400
rect 213360 0 213416 400
rect 214256 0 214312 400
rect 215152 0 215208 400
rect 216048 0 216104 400
rect 216944 0 217000 400
rect 217840 0 217896 400
rect 218736 0 218792 400
rect 219632 0 219688 400
rect 220528 0 220584 400
rect 221424 0 221480 400
rect 222320 0 222376 400
rect 223216 0 223272 400
rect 224112 0 224168 400
rect 225008 0 225064 400
rect 225904 0 225960 400
rect 226800 0 226856 400
rect 227696 0 227752 400
rect 228592 0 228648 400
rect 229488 0 229544 400
rect 230384 0 230440 400
rect 231280 0 231336 400
rect 232176 0 232232 400
rect 233072 0 233128 400
rect 233968 0 234024 400
rect 234864 0 234920 400
rect 235760 0 235816 400
rect 236656 0 236712 400
rect 237552 0 237608 400
rect 238448 0 238504 400
rect 239344 0 239400 400
rect 240240 0 240296 400
rect 241136 0 241192 400
rect 242032 0 242088 400
rect 242928 0 242984 400
rect 243824 0 243880 400
rect 244720 0 244776 400
rect 245616 0 245672 400
rect 246512 0 246568 400
rect 247408 0 247464 400
rect 248304 0 248360 400
rect 249200 0 249256 400
rect 250096 0 250152 400
rect 250992 0 251048 400
rect 251888 0 251944 400
rect 252784 0 252840 400
rect 253680 0 253736 400
rect 254576 0 254632 400
rect 255472 0 255528 400
rect 256368 0 256424 400
rect 257264 0 257320 400
rect 258160 0 258216 400
rect 259056 0 259112 400
rect 259952 0 260008 400
rect 260848 0 260904 400
rect 261744 0 261800 400
rect 262640 0 262696 400
rect 263536 0 263592 400
rect 264432 0 264488 400
rect 265328 0 265384 400
rect 266224 0 266280 400
rect 267120 0 267176 400
rect 268016 0 268072 400
rect 268912 0 268968 400
rect 269808 0 269864 400
rect 270704 0 270760 400
rect 271600 0 271656 400
rect 272496 0 272552 400
rect 273392 0 273448 400
rect 274288 0 274344 400
<< obsm2 >>
rect 966 430 278922 248155
rect 966 289 5458 430
rect 5574 289 6354 430
rect 6470 289 7250 430
rect 7366 289 8146 430
rect 8262 289 9042 430
rect 9158 289 9938 430
rect 10054 289 10834 430
rect 10950 289 11730 430
rect 11846 289 12626 430
rect 12742 289 13522 430
rect 13638 289 14418 430
rect 14534 289 15314 430
rect 15430 289 16210 430
rect 16326 289 17106 430
rect 17222 289 18002 430
rect 18118 289 18898 430
rect 19014 289 19794 430
rect 19910 289 20690 430
rect 20806 289 21586 430
rect 21702 289 22482 430
rect 22598 289 23378 430
rect 23494 289 24274 430
rect 24390 289 25170 430
rect 25286 289 26066 430
rect 26182 289 26962 430
rect 27078 289 27858 430
rect 27974 289 28754 430
rect 28870 289 29650 430
rect 29766 289 30546 430
rect 30662 289 31442 430
rect 31558 289 32338 430
rect 32454 289 33234 430
rect 33350 289 34130 430
rect 34246 289 35026 430
rect 35142 289 35922 430
rect 36038 289 36818 430
rect 36934 289 37714 430
rect 37830 289 38610 430
rect 38726 289 39506 430
rect 39622 289 40402 430
rect 40518 289 41298 430
rect 41414 289 42194 430
rect 42310 289 43090 430
rect 43206 289 43986 430
rect 44102 289 44882 430
rect 44998 289 45778 430
rect 45894 289 46674 430
rect 46790 289 47570 430
rect 47686 289 48466 430
rect 48582 289 49362 430
rect 49478 289 50258 430
rect 50374 289 51154 430
rect 51270 289 52050 430
rect 52166 289 52946 430
rect 53062 289 53842 430
rect 53958 289 54738 430
rect 54854 289 55634 430
rect 55750 289 56530 430
rect 56646 289 57426 430
rect 57542 289 58322 430
rect 58438 289 59218 430
rect 59334 289 60114 430
rect 60230 289 61010 430
rect 61126 289 61906 430
rect 62022 289 62802 430
rect 62918 289 63698 430
rect 63814 289 64594 430
rect 64710 289 65490 430
rect 65606 289 66386 430
rect 66502 289 67282 430
rect 67398 289 68178 430
rect 68294 289 69074 430
rect 69190 289 69970 430
rect 70086 289 70866 430
rect 70982 289 71762 430
rect 71878 289 72658 430
rect 72774 289 73554 430
rect 73670 289 74450 430
rect 74566 289 75346 430
rect 75462 289 76242 430
rect 76358 289 77138 430
rect 77254 289 78034 430
rect 78150 289 78930 430
rect 79046 289 79826 430
rect 79942 289 80722 430
rect 80838 289 81618 430
rect 81734 289 82514 430
rect 82630 289 83410 430
rect 83526 289 84306 430
rect 84422 289 85202 430
rect 85318 289 86098 430
rect 86214 289 86994 430
rect 87110 289 87890 430
rect 88006 289 88786 430
rect 88902 289 89682 430
rect 89798 289 90578 430
rect 90694 289 91474 430
rect 91590 289 92370 430
rect 92486 289 93266 430
rect 93382 289 94162 430
rect 94278 289 95058 430
rect 95174 289 95954 430
rect 96070 289 96850 430
rect 96966 289 97746 430
rect 97862 289 98642 430
rect 98758 289 99538 430
rect 99654 289 100434 430
rect 100550 289 101330 430
rect 101446 289 102226 430
rect 102342 289 103122 430
rect 103238 289 104018 430
rect 104134 289 104914 430
rect 105030 289 105810 430
rect 105926 289 106706 430
rect 106822 289 107602 430
rect 107718 289 108498 430
rect 108614 289 109394 430
rect 109510 289 110290 430
rect 110406 289 111186 430
rect 111302 289 112082 430
rect 112198 289 112978 430
rect 113094 289 113874 430
rect 113990 289 114770 430
rect 114886 289 115666 430
rect 115782 289 116562 430
rect 116678 289 117458 430
rect 117574 289 118354 430
rect 118470 289 119250 430
rect 119366 289 120146 430
rect 120262 289 121042 430
rect 121158 289 121938 430
rect 122054 289 122834 430
rect 122950 289 123730 430
rect 123846 289 124626 430
rect 124742 289 125522 430
rect 125638 289 126418 430
rect 126534 289 127314 430
rect 127430 289 128210 430
rect 128326 289 129106 430
rect 129222 289 130002 430
rect 130118 289 130898 430
rect 131014 289 131794 430
rect 131910 289 132690 430
rect 132806 289 133586 430
rect 133702 289 134482 430
rect 134598 289 135378 430
rect 135494 289 136274 430
rect 136390 289 137170 430
rect 137286 289 138066 430
rect 138182 289 138962 430
rect 139078 289 139858 430
rect 139974 289 140754 430
rect 140870 289 141650 430
rect 141766 289 142546 430
rect 142662 289 143442 430
rect 143558 289 144338 430
rect 144454 289 145234 430
rect 145350 289 146130 430
rect 146246 289 147026 430
rect 147142 289 147922 430
rect 148038 289 148818 430
rect 148934 289 149714 430
rect 149830 289 150610 430
rect 150726 289 151506 430
rect 151622 289 152402 430
rect 152518 289 153298 430
rect 153414 289 154194 430
rect 154310 289 155090 430
rect 155206 289 155986 430
rect 156102 289 156882 430
rect 156998 289 157778 430
rect 157894 289 158674 430
rect 158790 289 159570 430
rect 159686 289 160466 430
rect 160582 289 161362 430
rect 161478 289 162258 430
rect 162374 289 163154 430
rect 163270 289 164050 430
rect 164166 289 164946 430
rect 165062 289 165842 430
rect 165958 289 166738 430
rect 166854 289 167634 430
rect 167750 289 168530 430
rect 168646 289 169426 430
rect 169542 289 170322 430
rect 170438 289 171218 430
rect 171334 289 172114 430
rect 172230 289 173010 430
rect 173126 289 173906 430
rect 174022 289 174802 430
rect 174918 289 175698 430
rect 175814 289 176594 430
rect 176710 289 177490 430
rect 177606 289 178386 430
rect 178502 289 179282 430
rect 179398 289 180178 430
rect 180294 289 181074 430
rect 181190 289 181970 430
rect 182086 289 182866 430
rect 182982 289 183762 430
rect 183878 289 184658 430
rect 184774 289 185554 430
rect 185670 289 186450 430
rect 186566 289 187346 430
rect 187462 289 188242 430
rect 188358 289 189138 430
rect 189254 289 190034 430
rect 190150 289 190930 430
rect 191046 289 191826 430
rect 191942 289 192722 430
rect 192838 289 193618 430
rect 193734 289 194514 430
rect 194630 289 195410 430
rect 195526 289 196306 430
rect 196422 289 197202 430
rect 197318 289 198098 430
rect 198214 289 198994 430
rect 199110 289 199890 430
rect 200006 289 200786 430
rect 200902 289 201682 430
rect 201798 289 202578 430
rect 202694 289 203474 430
rect 203590 289 204370 430
rect 204486 289 205266 430
rect 205382 289 206162 430
rect 206278 289 207058 430
rect 207174 289 207954 430
rect 208070 289 208850 430
rect 208966 289 209746 430
rect 209862 289 210642 430
rect 210758 289 211538 430
rect 211654 289 212434 430
rect 212550 289 213330 430
rect 213446 289 214226 430
rect 214342 289 215122 430
rect 215238 289 216018 430
rect 216134 289 216914 430
rect 217030 289 217810 430
rect 217926 289 218706 430
rect 218822 289 219602 430
rect 219718 289 220498 430
rect 220614 289 221394 430
rect 221510 289 222290 430
rect 222406 289 223186 430
rect 223302 289 224082 430
rect 224198 289 224978 430
rect 225094 289 225874 430
rect 225990 289 226770 430
rect 226886 289 227666 430
rect 227782 289 228562 430
rect 228678 289 229458 430
rect 229574 289 230354 430
rect 230470 289 231250 430
rect 231366 289 232146 430
rect 232262 289 233042 430
rect 233158 289 233938 430
rect 234054 289 234834 430
rect 234950 289 235730 430
rect 235846 289 236626 430
rect 236742 289 237522 430
rect 237638 289 238418 430
rect 238534 289 239314 430
rect 239430 289 240210 430
rect 240326 289 241106 430
rect 241222 289 242002 430
rect 242118 289 242898 430
rect 243014 289 243794 430
rect 243910 289 244690 430
rect 244806 289 245586 430
rect 245702 289 246482 430
rect 246598 289 247378 430
rect 247494 289 248274 430
rect 248390 289 249170 430
rect 249286 289 250066 430
rect 250182 289 250962 430
rect 251078 289 251858 430
rect 251974 289 252754 430
rect 252870 289 253650 430
rect 253766 289 254546 430
rect 254662 289 255442 430
rect 255558 289 256338 430
rect 256454 289 257234 430
rect 257350 289 258130 430
rect 258246 289 259026 430
rect 259142 289 259922 430
rect 260038 289 260818 430
rect 260934 289 261714 430
rect 261830 289 262610 430
rect 262726 289 263506 430
rect 263622 289 264402 430
rect 264518 289 265298 430
rect 265414 289 266194 430
rect 266310 289 267090 430
rect 267206 289 267986 430
rect 268102 289 268882 430
rect 268998 289 269778 430
rect 269894 289 270674 430
rect 270790 289 271570 430
rect 271686 289 272466 430
rect 272582 289 273362 430
rect 273478 289 274258 430
rect 274374 289 278922 430
<< metal3 >>
rect 0 244720 400 244776
rect 279600 244720 280000 244776
rect 0 234304 400 234360
rect 279600 234304 280000 234360
rect 0 223888 400 223944
rect 279600 223888 280000 223944
rect 0 213472 400 213528
rect 279600 213472 280000 213528
rect 0 203056 400 203112
rect 279600 203056 280000 203112
rect 0 192640 400 192696
rect 279600 192640 280000 192696
rect 0 182224 400 182280
rect 279600 182224 280000 182280
rect 0 171808 400 171864
rect 279600 171808 280000 171864
rect 0 161392 400 161448
rect 279600 161392 280000 161448
rect 0 150976 400 151032
rect 279600 150976 280000 151032
rect 0 140560 400 140616
rect 279600 140560 280000 140616
rect 0 130144 400 130200
rect 279600 130144 280000 130200
rect 0 119728 400 119784
rect 279600 119728 280000 119784
rect 0 109312 400 109368
rect 279600 109312 280000 109368
rect 0 98896 400 98952
rect 279600 98896 280000 98952
rect 0 88480 400 88536
rect 279600 88480 280000 88536
rect 0 78064 400 78120
rect 279600 78064 280000 78120
rect 0 67648 400 67704
rect 279600 67648 280000 67704
rect 0 57232 400 57288
rect 279600 57232 280000 57288
rect 0 46816 400 46872
rect 279600 46816 280000 46872
rect 0 36400 400 36456
rect 279600 36400 280000 36456
rect 0 25984 400 26040
rect 279600 25984 280000 26040
rect 0 15568 400 15624
rect 279600 15568 280000 15624
rect 0 5152 400 5208
rect 279600 5152 280000 5208
<< obsm3 >>
rect 400 244806 279650 248150
rect 430 244690 279570 244806
rect 400 234390 279650 244690
rect 430 234274 279570 234390
rect 400 223974 279650 234274
rect 430 223858 279570 223974
rect 400 213558 279650 223858
rect 430 213442 279570 213558
rect 400 203142 279650 213442
rect 430 203026 279570 203142
rect 400 192726 279650 203026
rect 430 192610 279570 192726
rect 400 182310 279650 192610
rect 430 182194 279570 182310
rect 400 171894 279650 182194
rect 430 171778 279570 171894
rect 400 161478 279650 171778
rect 430 161362 279570 161478
rect 400 151062 279650 161362
rect 430 150946 279570 151062
rect 400 140646 279650 150946
rect 430 140530 279570 140646
rect 400 130230 279650 140530
rect 430 130114 279570 130230
rect 400 119814 279650 130114
rect 430 119698 279570 119814
rect 400 109398 279650 119698
rect 430 109282 279570 109398
rect 400 98982 279650 109282
rect 430 98866 279570 98982
rect 400 88566 279650 98866
rect 430 88450 279570 88566
rect 400 78150 279650 88450
rect 430 78034 279570 78150
rect 400 67734 279650 78034
rect 430 67618 279570 67734
rect 400 57318 279650 67618
rect 430 57202 279570 57318
rect 400 46902 279650 57202
rect 430 46786 279570 46902
rect 400 36486 279650 46786
rect 430 36370 279570 36486
rect 400 26070 279650 36370
rect 430 25954 279570 26070
rect 400 15654 279650 25954
rect 430 15538 279570 15654
rect 400 5238 279650 15538
rect 430 5122 279570 5238
rect 400 294 279650 5122
<< metal4 >>
rect 2224 1538 2384 248166
rect 9904 1538 10064 248166
rect 17584 1538 17744 248166
rect 25264 1538 25424 248166
rect 32944 1538 33104 248166
rect 40624 1538 40784 248166
rect 48304 1538 48464 248166
rect 55984 1538 56144 248166
rect 63664 1538 63824 248166
rect 71344 1538 71504 248166
rect 79024 1538 79184 248166
rect 86704 1538 86864 248166
rect 94384 1538 94544 248166
rect 102064 1538 102224 248166
rect 109744 1538 109904 248166
rect 117424 1538 117584 248166
rect 125104 1538 125264 248166
rect 132784 1538 132944 248166
rect 140464 1538 140624 248166
rect 148144 1538 148304 248166
rect 155824 1538 155984 248166
rect 163504 1538 163664 248166
rect 171184 1538 171344 248166
rect 178864 1538 179024 248166
rect 186544 1538 186704 248166
rect 194224 1538 194384 248166
rect 201904 1538 202064 248166
rect 209584 1538 209744 248166
rect 217264 1538 217424 248166
rect 224944 1538 225104 248166
rect 232624 1538 232784 248166
rect 240304 1538 240464 248166
rect 247984 1538 248144 248166
rect 255664 1538 255824 248166
rect 263344 1538 263504 248166
rect 271024 1538 271184 248166
rect 278704 1538 278864 248166
<< obsm4 >>
rect 126238 1508 132754 8559
rect 132974 1508 140434 8559
rect 140654 1508 146986 8559
rect 126238 345 146986 1508
<< labels >>
rlabel metal3 s 279600 5152 280000 5208 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 182224 400 182280 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 150976 400 151032 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 119728 400 119784 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 0 88480 400 88536 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 0 57232 400 57288 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 25984 400 26040 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 279600 36400 280000 36456 6 io_in[1]
port 8 nsew signal input
rlabel metal3 s 279600 67648 280000 67704 6 io_in[2]
port 9 nsew signal input
rlabel metal3 s 279600 98896 280000 98952 6 io_in[3]
port 10 nsew signal input
rlabel metal3 s 279600 130144 280000 130200 6 io_in[4]
port 11 nsew signal input
rlabel metal3 s 279600 161392 280000 161448 6 io_in[5]
port 12 nsew signal input
rlabel metal3 s 279600 192640 280000 192696 6 io_in[6]
port 13 nsew signal input
rlabel metal3 s 279600 223888 280000 223944 6 io_in[7]
port 14 nsew signal input
rlabel metal3 s 0 244720 400 244776 6 io_in[8]
port 15 nsew signal input
rlabel metal3 s 0 213472 400 213528 6 io_in[9]
port 16 nsew signal input
rlabel metal3 s 279600 25984 280000 26040 6 io_oeb[0]
port 17 nsew signal output
rlabel metal3 s 0 161392 400 161448 6 io_oeb[10]
port 18 nsew signal output
rlabel metal3 s 0 130144 400 130200 6 io_oeb[11]
port 19 nsew signal output
rlabel metal3 s 0 98896 400 98952 6 io_oeb[12]
port 20 nsew signal output
rlabel metal3 s 0 67648 400 67704 6 io_oeb[13]
port 21 nsew signal output
rlabel metal3 s 0 36400 400 36456 6 io_oeb[14]
port 22 nsew signal output
rlabel metal3 s 0 5152 400 5208 6 io_oeb[15]
port 23 nsew signal output
rlabel metal3 s 279600 57232 280000 57288 6 io_oeb[1]
port 24 nsew signal output
rlabel metal3 s 279600 88480 280000 88536 6 io_oeb[2]
port 25 nsew signal output
rlabel metal3 s 279600 119728 280000 119784 6 io_oeb[3]
port 26 nsew signal output
rlabel metal3 s 279600 150976 280000 151032 6 io_oeb[4]
port 27 nsew signal output
rlabel metal3 s 279600 182224 280000 182280 6 io_oeb[5]
port 28 nsew signal output
rlabel metal3 s 279600 213472 280000 213528 6 io_oeb[6]
port 29 nsew signal output
rlabel metal3 s 279600 244720 280000 244776 6 io_oeb[7]
port 30 nsew signal output
rlabel metal3 s 0 223888 400 223944 6 io_oeb[8]
port 31 nsew signal output
rlabel metal3 s 0 192640 400 192696 6 io_oeb[9]
port 32 nsew signal output
rlabel metal3 s 279600 15568 280000 15624 6 io_out[0]
port 33 nsew signal output
rlabel metal3 s 0 171808 400 171864 6 io_out[10]
port 34 nsew signal output
rlabel metal3 s 0 140560 400 140616 6 io_out[11]
port 35 nsew signal output
rlabel metal3 s 0 109312 400 109368 6 io_out[12]
port 36 nsew signal output
rlabel metal3 s 0 78064 400 78120 6 io_out[13]
port 37 nsew signal output
rlabel metal3 s 0 46816 400 46872 6 io_out[14]
port 38 nsew signal output
rlabel metal3 s 0 15568 400 15624 6 io_out[15]
port 39 nsew signal output
rlabel metal3 s 279600 46816 280000 46872 6 io_out[1]
port 40 nsew signal output
rlabel metal3 s 279600 78064 280000 78120 6 io_out[2]
port 41 nsew signal output
rlabel metal3 s 279600 109312 280000 109368 6 io_out[3]
port 42 nsew signal output
rlabel metal3 s 279600 140560 280000 140616 6 io_out[4]
port 43 nsew signal output
rlabel metal3 s 279600 171808 280000 171864 6 io_out[5]
port 44 nsew signal output
rlabel metal3 s 279600 203056 280000 203112 6 io_out[6]
port 45 nsew signal output
rlabel metal3 s 279600 234304 280000 234360 6 io_out[7]
port 46 nsew signal output
rlabel metal3 s 0 234304 400 234360 6 io_out[8]
port 47 nsew signal output
rlabel metal3 s 0 203056 400 203112 6 io_out[9]
port 48 nsew signal output
rlabel metal2 s 272496 0 272552 400 6 irq[0]
port 49 nsew signal output
rlabel metal2 s 273392 0 273448 400 6 irq[1]
port 50 nsew signal output
rlabel metal2 s 274288 0 274344 400 6 irq[2]
port 51 nsew signal output
rlabel metal2 s 100464 0 100520 400 6 la_data_in[0]
port 52 nsew signal input
rlabel metal2 s 127344 0 127400 400 6 la_data_in[10]
port 53 nsew signal input
rlabel metal2 s 130032 0 130088 400 6 la_data_in[11]
port 54 nsew signal input
rlabel metal2 s 132720 0 132776 400 6 la_data_in[12]
port 55 nsew signal input
rlabel metal2 s 135408 0 135464 400 6 la_data_in[13]
port 56 nsew signal input
rlabel metal2 s 138096 0 138152 400 6 la_data_in[14]
port 57 nsew signal input
rlabel metal2 s 140784 0 140840 400 6 la_data_in[15]
port 58 nsew signal input
rlabel metal2 s 143472 0 143528 400 6 la_data_in[16]
port 59 nsew signal input
rlabel metal2 s 146160 0 146216 400 6 la_data_in[17]
port 60 nsew signal input
rlabel metal2 s 148848 0 148904 400 6 la_data_in[18]
port 61 nsew signal input
rlabel metal2 s 151536 0 151592 400 6 la_data_in[19]
port 62 nsew signal input
rlabel metal2 s 103152 0 103208 400 6 la_data_in[1]
port 63 nsew signal input
rlabel metal2 s 154224 0 154280 400 6 la_data_in[20]
port 64 nsew signal input
rlabel metal2 s 156912 0 156968 400 6 la_data_in[21]
port 65 nsew signal input
rlabel metal2 s 159600 0 159656 400 6 la_data_in[22]
port 66 nsew signal input
rlabel metal2 s 162288 0 162344 400 6 la_data_in[23]
port 67 nsew signal input
rlabel metal2 s 164976 0 165032 400 6 la_data_in[24]
port 68 nsew signal input
rlabel metal2 s 167664 0 167720 400 6 la_data_in[25]
port 69 nsew signal input
rlabel metal2 s 170352 0 170408 400 6 la_data_in[26]
port 70 nsew signal input
rlabel metal2 s 173040 0 173096 400 6 la_data_in[27]
port 71 nsew signal input
rlabel metal2 s 175728 0 175784 400 6 la_data_in[28]
port 72 nsew signal input
rlabel metal2 s 178416 0 178472 400 6 la_data_in[29]
port 73 nsew signal input
rlabel metal2 s 105840 0 105896 400 6 la_data_in[2]
port 74 nsew signal input
rlabel metal2 s 181104 0 181160 400 6 la_data_in[30]
port 75 nsew signal input
rlabel metal2 s 183792 0 183848 400 6 la_data_in[31]
port 76 nsew signal input
rlabel metal2 s 186480 0 186536 400 6 la_data_in[32]
port 77 nsew signal input
rlabel metal2 s 189168 0 189224 400 6 la_data_in[33]
port 78 nsew signal input
rlabel metal2 s 191856 0 191912 400 6 la_data_in[34]
port 79 nsew signal input
rlabel metal2 s 194544 0 194600 400 6 la_data_in[35]
port 80 nsew signal input
rlabel metal2 s 197232 0 197288 400 6 la_data_in[36]
port 81 nsew signal input
rlabel metal2 s 199920 0 199976 400 6 la_data_in[37]
port 82 nsew signal input
rlabel metal2 s 202608 0 202664 400 6 la_data_in[38]
port 83 nsew signal input
rlabel metal2 s 205296 0 205352 400 6 la_data_in[39]
port 84 nsew signal input
rlabel metal2 s 108528 0 108584 400 6 la_data_in[3]
port 85 nsew signal input
rlabel metal2 s 207984 0 208040 400 6 la_data_in[40]
port 86 nsew signal input
rlabel metal2 s 210672 0 210728 400 6 la_data_in[41]
port 87 nsew signal input
rlabel metal2 s 213360 0 213416 400 6 la_data_in[42]
port 88 nsew signal input
rlabel metal2 s 216048 0 216104 400 6 la_data_in[43]
port 89 nsew signal input
rlabel metal2 s 218736 0 218792 400 6 la_data_in[44]
port 90 nsew signal input
rlabel metal2 s 221424 0 221480 400 6 la_data_in[45]
port 91 nsew signal input
rlabel metal2 s 224112 0 224168 400 6 la_data_in[46]
port 92 nsew signal input
rlabel metal2 s 226800 0 226856 400 6 la_data_in[47]
port 93 nsew signal input
rlabel metal2 s 229488 0 229544 400 6 la_data_in[48]
port 94 nsew signal input
rlabel metal2 s 232176 0 232232 400 6 la_data_in[49]
port 95 nsew signal input
rlabel metal2 s 111216 0 111272 400 6 la_data_in[4]
port 96 nsew signal input
rlabel metal2 s 234864 0 234920 400 6 la_data_in[50]
port 97 nsew signal input
rlabel metal2 s 237552 0 237608 400 6 la_data_in[51]
port 98 nsew signal input
rlabel metal2 s 240240 0 240296 400 6 la_data_in[52]
port 99 nsew signal input
rlabel metal2 s 242928 0 242984 400 6 la_data_in[53]
port 100 nsew signal input
rlabel metal2 s 245616 0 245672 400 6 la_data_in[54]
port 101 nsew signal input
rlabel metal2 s 248304 0 248360 400 6 la_data_in[55]
port 102 nsew signal input
rlabel metal2 s 250992 0 251048 400 6 la_data_in[56]
port 103 nsew signal input
rlabel metal2 s 253680 0 253736 400 6 la_data_in[57]
port 104 nsew signal input
rlabel metal2 s 256368 0 256424 400 6 la_data_in[58]
port 105 nsew signal input
rlabel metal2 s 259056 0 259112 400 6 la_data_in[59]
port 106 nsew signal input
rlabel metal2 s 113904 0 113960 400 6 la_data_in[5]
port 107 nsew signal input
rlabel metal2 s 261744 0 261800 400 6 la_data_in[60]
port 108 nsew signal input
rlabel metal2 s 264432 0 264488 400 6 la_data_in[61]
port 109 nsew signal input
rlabel metal2 s 267120 0 267176 400 6 la_data_in[62]
port 110 nsew signal input
rlabel metal2 s 269808 0 269864 400 6 la_data_in[63]
port 111 nsew signal input
rlabel metal2 s 116592 0 116648 400 6 la_data_in[6]
port 112 nsew signal input
rlabel metal2 s 119280 0 119336 400 6 la_data_in[7]
port 113 nsew signal input
rlabel metal2 s 121968 0 122024 400 6 la_data_in[8]
port 114 nsew signal input
rlabel metal2 s 124656 0 124712 400 6 la_data_in[9]
port 115 nsew signal input
rlabel metal2 s 101360 0 101416 400 6 la_data_out[0]
port 116 nsew signal output
rlabel metal2 s 128240 0 128296 400 6 la_data_out[10]
port 117 nsew signal output
rlabel metal2 s 130928 0 130984 400 6 la_data_out[11]
port 118 nsew signal output
rlabel metal2 s 133616 0 133672 400 6 la_data_out[12]
port 119 nsew signal output
rlabel metal2 s 136304 0 136360 400 6 la_data_out[13]
port 120 nsew signal output
rlabel metal2 s 138992 0 139048 400 6 la_data_out[14]
port 121 nsew signal output
rlabel metal2 s 141680 0 141736 400 6 la_data_out[15]
port 122 nsew signal output
rlabel metal2 s 144368 0 144424 400 6 la_data_out[16]
port 123 nsew signal output
rlabel metal2 s 147056 0 147112 400 6 la_data_out[17]
port 124 nsew signal output
rlabel metal2 s 149744 0 149800 400 6 la_data_out[18]
port 125 nsew signal output
rlabel metal2 s 152432 0 152488 400 6 la_data_out[19]
port 126 nsew signal output
rlabel metal2 s 104048 0 104104 400 6 la_data_out[1]
port 127 nsew signal output
rlabel metal2 s 155120 0 155176 400 6 la_data_out[20]
port 128 nsew signal output
rlabel metal2 s 157808 0 157864 400 6 la_data_out[21]
port 129 nsew signal output
rlabel metal2 s 160496 0 160552 400 6 la_data_out[22]
port 130 nsew signal output
rlabel metal2 s 163184 0 163240 400 6 la_data_out[23]
port 131 nsew signal output
rlabel metal2 s 165872 0 165928 400 6 la_data_out[24]
port 132 nsew signal output
rlabel metal2 s 168560 0 168616 400 6 la_data_out[25]
port 133 nsew signal output
rlabel metal2 s 171248 0 171304 400 6 la_data_out[26]
port 134 nsew signal output
rlabel metal2 s 173936 0 173992 400 6 la_data_out[27]
port 135 nsew signal output
rlabel metal2 s 176624 0 176680 400 6 la_data_out[28]
port 136 nsew signal output
rlabel metal2 s 179312 0 179368 400 6 la_data_out[29]
port 137 nsew signal output
rlabel metal2 s 106736 0 106792 400 6 la_data_out[2]
port 138 nsew signal output
rlabel metal2 s 182000 0 182056 400 6 la_data_out[30]
port 139 nsew signal output
rlabel metal2 s 184688 0 184744 400 6 la_data_out[31]
port 140 nsew signal output
rlabel metal2 s 187376 0 187432 400 6 la_data_out[32]
port 141 nsew signal output
rlabel metal2 s 190064 0 190120 400 6 la_data_out[33]
port 142 nsew signal output
rlabel metal2 s 192752 0 192808 400 6 la_data_out[34]
port 143 nsew signal output
rlabel metal2 s 195440 0 195496 400 6 la_data_out[35]
port 144 nsew signal output
rlabel metal2 s 198128 0 198184 400 6 la_data_out[36]
port 145 nsew signal output
rlabel metal2 s 200816 0 200872 400 6 la_data_out[37]
port 146 nsew signal output
rlabel metal2 s 203504 0 203560 400 6 la_data_out[38]
port 147 nsew signal output
rlabel metal2 s 206192 0 206248 400 6 la_data_out[39]
port 148 nsew signal output
rlabel metal2 s 109424 0 109480 400 6 la_data_out[3]
port 149 nsew signal output
rlabel metal2 s 208880 0 208936 400 6 la_data_out[40]
port 150 nsew signal output
rlabel metal2 s 211568 0 211624 400 6 la_data_out[41]
port 151 nsew signal output
rlabel metal2 s 214256 0 214312 400 6 la_data_out[42]
port 152 nsew signal output
rlabel metal2 s 216944 0 217000 400 6 la_data_out[43]
port 153 nsew signal output
rlabel metal2 s 219632 0 219688 400 6 la_data_out[44]
port 154 nsew signal output
rlabel metal2 s 222320 0 222376 400 6 la_data_out[45]
port 155 nsew signal output
rlabel metal2 s 225008 0 225064 400 6 la_data_out[46]
port 156 nsew signal output
rlabel metal2 s 227696 0 227752 400 6 la_data_out[47]
port 157 nsew signal output
rlabel metal2 s 230384 0 230440 400 6 la_data_out[48]
port 158 nsew signal output
rlabel metal2 s 233072 0 233128 400 6 la_data_out[49]
port 159 nsew signal output
rlabel metal2 s 112112 0 112168 400 6 la_data_out[4]
port 160 nsew signal output
rlabel metal2 s 235760 0 235816 400 6 la_data_out[50]
port 161 nsew signal output
rlabel metal2 s 238448 0 238504 400 6 la_data_out[51]
port 162 nsew signal output
rlabel metal2 s 241136 0 241192 400 6 la_data_out[52]
port 163 nsew signal output
rlabel metal2 s 243824 0 243880 400 6 la_data_out[53]
port 164 nsew signal output
rlabel metal2 s 246512 0 246568 400 6 la_data_out[54]
port 165 nsew signal output
rlabel metal2 s 249200 0 249256 400 6 la_data_out[55]
port 166 nsew signal output
rlabel metal2 s 251888 0 251944 400 6 la_data_out[56]
port 167 nsew signal output
rlabel metal2 s 254576 0 254632 400 6 la_data_out[57]
port 168 nsew signal output
rlabel metal2 s 257264 0 257320 400 6 la_data_out[58]
port 169 nsew signal output
rlabel metal2 s 259952 0 260008 400 6 la_data_out[59]
port 170 nsew signal output
rlabel metal2 s 114800 0 114856 400 6 la_data_out[5]
port 171 nsew signal output
rlabel metal2 s 262640 0 262696 400 6 la_data_out[60]
port 172 nsew signal output
rlabel metal2 s 265328 0 265384 400 6 la_data_out[61]
port 173 nsew signal output
rlabel metal2 s 268016 0 268072 400 6 la_data_out[62]
port 174 nsew signal output
rlabel metal2 s 270704 0 270760 400 6 la_data_out[63]
port 175 nsew signal output
rlabel metal2 s 117488 0 117544 400 6 la_data_out[6]
port 176 nsew signal output
rlabel metal2 s 120176 0 120232 400 6 la_data_out[7]
port 177 nsew signal output
rlabel metal2 s 122864 0 122920 400 6 la_data_out[8]
port 178 nsew signal output
rlabel metal2 s 125552 0 125608 400 6 la_data_out[9]
port 179 nsew signal output
rlabel metal2 s 102256 0 102312 400 6 la_oenb[0]
port 180 nsew signal input
rlabel metal2 s 129136 0 129192 400 6 la_oenb[10]
port 181 nsew signal input
rlabel metal2 s 131824 0 131880 400 6 la_oenb[11]
port 182 nsew signal input
rlabel metal2 s 134512 0 134568 400 6 la_oenb[12]
port 183 nsew signal input
rlabel metal2 s 137200 0 137256 400 6 la_oenb[13]
port 184 nsew signal input
rlabel metal2 s 139888 0 139944 400 6 la_oenb[14]
port 185 nsew signal input
rlabel metal2 s 142576 0 142632 400 6 la_oenb[15]
port 186 nsew signal input
rlabel metal2 s 145264 0 145320 400 6 la_oenb[16]
port 187 nsew signal input
rlabel metal2 s 147952 0 148008 400 6 la_oenb[17]
port 188 nsew signal input
rlabel metal2 s 150640 0 150696 400 6 la_oenb[18]
port 189 nsew signal input
rlabel metal2 s 153328 0 153384 400 6 la_oenb[19]
port 190 nsew signal input
rlabel metal2 s 104944 0 105000 400 6 la_oenb[1]
port 191 nsew signal input
rlabel metal2 s 156016 0 156072 400 6 la_oenb[20]
port 192 nsew signal input
rlabel metal2 s 158704 0 158760 400 6 la_oenb[21]
port 193 nsew signal input
rlabel metal2 s 161392 0 161448 400 6 la_oenb[22]
port 194 nsew signal input
rlabel metal2 s 164080 0 164136 400 6 la_oenb[23]
port 195 nsew signal input
rlabel metal2 s 166768 0 166824 400 6 la_oenb[24]
port 196 nsew signal input
rlabel metal2 s 169456 0 169512 400 6 la_oenb[25]
port 197 nsew signal input
rlabel metal2 s 172144 0 172200 400 6 la_oenb[26]
port 198 nsew signal input
rlabel metal2 s 174832 0 174888 400 6 la_oenb[27]
port 199 nsew signal input
rlabel metal2 s 177520 0 177576 400 6 la_oenb[28]
port 200 nsew signal input
rlabel metal2 s 180208 0 180264 400 6 la_oenb[29]
port 201 nsew signal input
rlabel metal2 s 107632 0 107688 400 6 la_oenb[2]
port 202 nsew signal input
rlabel metal2 s 182896 0 182952 400 6 la_oenb[30]
port 203 nsew signal input
rlabel metal2 s 185584 0 185640 400 6 la_oenb[31]
port 204 nsew signal input
rlabel metal2 s 188272 0 188328 400 6 la_oenb[32]
port 205 nsew signal input
rlabel metal2 s 190960 0 191016 400 6 la_oenb[33]
port 206 nsew signal input
rlabel metal2 s 193648 0 193704 400 6 la_oenb[34]
port 207 nsew signal input
rlabel metal2 s 196336 0 196392 400 6 la_oenb[35]
port 208 nsew signal input
rlabel metal2 s 199024 0 199080 400 6 la_oenb[36]
port 209 nsew signal input
rlabel metal2 s 201712 0 201768 400 6 la_oenb[37]
port 210 nsew signal input
rlabel metal2 s 204400 0 204456 400 6 la_oenb[38]
port 211 nsew signal input
rlabel metal2 s 207088 0 207144 400 6 la_oenb[39]
port 212 nsew signal input
rlabel metal2 s 110320 0 110376 400 6 la_oenb[3]
port 213 nsew signal input
rlabel metal2 s 209776 0 209832 400 6 la_oenb[40]
port 214 nsew signal input
rlabel metal2 s 212464 0 212520 400 6 la_oenb[41]
port 215 nsew signal input
rlabel metal2 s 215152 0 215208 400 6 la_oenb[42]
port 216 nsew signal input
rlabel metal2 s 217840 0 217896 400 6 la_oenb[43]
port 217 nsew signal input
rlabel metal2 s 220528 0 220584 400 6 la_oenb[44]
port 218 nsew signal input
rlabel metal2 s 223216 0 223272 400 6 la_oenb[45]
port 219 nsew signal input
rlabel metal2 s 225904 0 225960 400 6 la_oenb[46]
port 220 nsew signal input
rlabel metal2 s 228592 0 228648 400 6 la_oenb[47]
port 221 nsew signal input
rlabel metal2 s 231280 0 231336 400 6 la_oenb[48]
port 222 nsew signal input
rlabel metal2 s 233968 0 234024 400 6 la_oenb[49]
port 223 nsew signal input
rlabel metal2 s 113008 0 113064 400 6 la_oenb[4]
port 224 nsew signal input
rlabel metal2 s 236656 0 236712 400 6 la_oenb[50]
port 225 nsew signal input
rlabel metal2 s 239344 0 239400 400 6 la_oenb[51]
port 226 nsew signal input
rlabel metal2 s 242032 0 242088 400 6 la_oenb[52]
port 227 nsew signal input
rlabel metal2 s 244720 0 244776 400 6 la_oenb[53]
port 228 nsew signal input
rlabel metal2 s 247408 0 247464 400 6 la_oenb[54]
port 229 nsew signal input
rlabel metal2 s 250096 0 250152 400 6 la_oenb[55]
port 230 nsew signal input
rlabel metal2 s 252784 0 252840 400 6 la_oenb[56]
port 231 nsew signal input
rlabel metal2 s 255472 0 255528 400 6 la_oenb[57]
port 232 nsew signal input
rlabel metal2 s 258160 0 258216 400 6 la_oenb[58]
port 233 nsew signal input
rlabel metal2 s 260848 0 260904 400 6 la_oenb[59]
port 234 nsew signal input
rlabel metal2 s 115696 0 115752 400 6 la_oenb[5]
port 235 nsew signal input
rlabel metal2 s 263536 0 263592 400 6 la_oenb[60]
port 236 nsew signal input
rlabel metal2 s 266224 0 266280 400 6 la_oenb[61]
port 237 nsew signal input
rlabel metal2 s 268912 0 268968 400 6 la_oenb[62]
port 238 nsew signal input
rlabel metal2 s 271600 0 271656 400 6 la_oenb[63]
port 239 nsew signal input
rlabel metal2 s 118384 0 118440 400 6 la_oenb[6]
port 240 nsew signal input
rlabel metal2 s 121072 0 121128 400 6 la_oenb[7]
port 241 nsew signal input
rlabel metal2 s 123760 0 123816 400 6 la_oenb[8]
port 242 nsew signal input
rlabel metal2 s 126448 0 126504 400 6 la_oenb[9]
port 243 nsew signal input
rlabel metal4 s 2224 1538 2384 248166 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 248166 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 248166 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 248166 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 248166 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 248166 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 248166 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 248166 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 248166 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 248166 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 248166 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 248166 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 248166 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 248166 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 248166 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 248166 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 248166 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 263344 1538 263504 248166 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 278704 1538 278864 248166 6 vdd
port 244 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 248166 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 248166 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 248166 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 248166 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 248166 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 248166 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 248166 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 248166 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 248166 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 248166 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 248166 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 248166 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 248166 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 248166 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 248166 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 248166 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 255664 1538 255824 248166 6 vss
port 245 nsew ground bidirectional
rlabel metal4 s 271024 1538 271184 248166 6 vss
port 245 nsew ground bidirectional
rlabel metal2 s 5488 0 5544 400 6 wb_clk_i
port 246 nsew signal input
rlabel metal2 s 6384 0 6440 400 6 wb_rst_i
port 247 nsew signal input
rlabel metal2 s 7280 0 7336 400 6 wbs_ack_o
port 248 nsew signal output
rlabel metal2 s 10864 0 10920 400 6 wbs_adr_i[0]
port 249 nsew signal input
rlabel metal2 s 41328 0 41384 400 6 wbs_adr_i[10]
port 250 nsew signal input
rlabel metal2 s 44016 0 44072 400 6 wbs_adr_i[11]
port 251 nsew signal input
rlabel metal2 s 46704 0 46760 400 6 wbs_adr_i[12]
port 252 nsew signal input
rlabel metal2 s 49392 0 49448 400 6 wbs_adr_i[13]
port 253 nsew signal input
rlabel metal2 s 52080 0 52136 400 6 wbs_adr_i[14]
port 254 nsew signal input
rlabel metal2 s 54768 0 54824 400 6 wbs_adr_i[15]
port 255 nsew signal input
rlabel metal2 s 57456 0 57512 400 6 wbs_adr_i[16]
port 256 nsew signal input
rlabel metal2 s 60144 0 60200 400 6 wbs_adr_i[17]
port 257 nsew signal input
rlabel metal2 s 62832 0 62888 400 6 wbs_adr_i[18]
port 258 nsew signal input
rlabel metal2 s 65520 0 65576 400 6 wbs_adr_i[19]
port 259 nsew signal input
rlabel metal2 s 14448 0 14504 400 6 wbs_adr_i[1]
port 260 nsew signal input
rlabel metal2 s 68208 0 68264 400 6 wbs_adr_i[20]
port 261 nsew signal input
rlabel metal2 s 70896 0 70952 400 6 wbs_adr_i[21]
port 262 nsew signal input
rlabel metal2 s 73584 0 73640 400 6 wbs_adr_i[22]
port 263 nsew signal input
rlabel metal2 s 76272 0 76328 400 6 wbs_adr_i[23]
port 264 nsew signal input
rlabel metal2 s 78960 0 79016 400 6 wbs_adr_i[24]
port 265 nsew signal input
rlabel metal2 s 81648 0 81704 400 6 wbs_adr_i[25]
port 266 nsew signal input
rlabel metal2 s 84336 0 84392 400 6 wbs_adr_i[26]
port 267 nsew signal input
rlabel metal2 s 87024 0 87080 400 6 wbs_adr_i[27]
port 268 nsew signal input
rlabel metal2 s 89712 0 89768 400 6 wbs_adr_i[28]
port 269 nsew signal input
rlabel metal2 s 92400 0 92456 400 6 wbs_adr_i[29]
port 270 nsew signal input
rlabel metal2 s 18032 0 18088 400 6 wbs_adr_i[2]
port 271 nsew signal input
rlabel metal2 s 95088 0 95144 400 6 wbs_adr_i[30]
port 272 nsew signal input
rlabel metal2 s 97776 0 97832 400 6 wbs_adr_i[31]
port 273 nsew signal input
rlabel metal2 s 21616 0 21672 400 6 wbs_adr_i[3]
port 274 nsew signal input
rlabel metal2 s 25200 0 25256 400 6 wbs_adr_i[4]
port 275 nsew signal input
rlabel metal2 s 27888 0 27944 400 6 wbs_adr_i[5]
port 276 nsew signal input
rlabel metal2 s 30576 0 30632 400 6 wbs_adr_i[6]
port 277 nsew signal input
rlabel metal2 s 33264 0 33320 400 6 wbs_adr_i[7]
port 278 nsew signal input
rlabel metal2 s 35952 0 36008 400 6 wbs_adr_i[8]
port 279 nsew signal input
rlabel metal2 s 38640 0 38696 400 6 wbs_adr_i[9]
port 280 nsew signal input
rlabel metal2 s 8176 0 8232 400 6 wbs_cyc_i
port 281 nsew signal input
rlabel metal2 s 11760 0 11816 400 6 wbs_dat_i[0]
port 282 nsew signal input
rlabel metal2 s 42224 0 42280 400 6 wbs_dat_i[10]
port 283 nsew signal input
rlabel metal2 s 44912 0 44968 400 6 wbs_dat_i[11]
port 284 nsew signal input
rlabel metal2 s 47600 0 47656 400 6 wbs_dat_i[12]
port 285 nsew signal input
rlabel metal2 s 50288 0 50344 400 6 wbs_dat_i[13]
port 286 nsew signal input
rlabel metal2 s 52976 0 53032 400 6 wbs_dat_i[14]
port 287 nsew signal input
rlabel metal2 s 55664 0 55720 400 6 wbs_dat_i[15]
port 288 nsew signal input
rlabel metal2 s 58352 0 58408 400 6 wbs_dat_i[16]
port 289 nsew signal input
rlabel metal2 s 61040 0 61096 400 6 wbs_dat_i[17]
port 290 nsew signal input
rlabel metal2 s 63728 0 63784 400 6 wbs_dat_i[18]
port 291 nsew signal input
rlabel metal2 s 66416 0 66472 400 6 wbs_dat_i[19]
port 292 nsew signal input
rlabel metal2 s 15344 0 15400 400 6 wbs_dat_i[1]
port 293 nsew signal input
rlabel metal2 s 69104 0 69160 400 6 wbs_dat_i[20]
port 294 nsew signal input
rlabel metal2 s 71792 0 71848 400 6 wbs_dat_i[21]
port 295 nsew signal input
rlabel metal2 s 74480 0 74536 400 6 wbs_dat_i[22]
port 296 nsew signal input
rlabel metal2 s 77168 0 77224 400 6 wbs_dat_i[23]
port 297 nsew signal input
rlabel metal2 s 79856 0 79912 400 6 wbs_dat_i[24]
port 298 nsew signal input
rlabel metal2 s 82544 0 82600 400 6 wbs_dat_i[25]
port 299 nsew signal input
rlabel metal2 s 85232 0 85288 400 6 wbs_dat_i[26]
port 300 nsew signal input
rlabel metal2 s 87920 0 87976 400 6 wbs_dat_i[27]
port 301 nsew signal input
rlabel metal2 s 90608 0 90664 400 6 wbs_dat_i[28]
port 302 nsew signal input
rlabel metal2 s 93296 0 93352 400 6 wbs_dat_i[29]
port 303 nsew signal input
rlabel metal2 s 18928 0 18984 400 6 wbs_dat_i[2]
port 304 nsew signal input
rlabel metal2 s 95984 0 96040 400 6 wbs_dat_i[30]
port 305 nsew signal input
rlabel metal2 s 98672 0 98728 400 6 wbs_dat_i[31]
port 306 nsew signal input
rlabel metal2 s 22512 0 22568 400 6 wbs_dat_i[3]
port 307 nsew signal input
rlabel metal2 s 26096 0 26152 400 6 wbs_dat_i[4]
port 308 nsew signal input
rlabel metal2 s 28784 0 28840 400 6 wbs_dat_i[5]
port 309 nsew signal input
rlabel metal2 s 31472 0 31528 400 6 wbs_dat_i[6]
port 310 nsew signal input
rlabel metal2 s 34160 0 34216 400 6 wbs_dat_i[7]
port 311 nsew signal input
rlabel metal2 s 36848 0 36904 400 6 wbs_dat_i[8]
port 312 nsew signal input
rlabel metal2 s 39536 0 39592 400 6 wbs_dat_i[9]
port 313 nsew signal input
rlabel metal2 s 12656 0 12712 400 6 wbs_dat_o[0]
port 314 nsew signal output
rlabel metal2 s 43120 0 43176 400 6 wbs_dat_o[10]
port 315 nsew signal output
rlabel metal2 s 45808 0 45864 400 6 wbs_dat_o[11]
port 316 nsew signal output
rlabel metal2 s 48496 0 48552 400 6 wbs_dat_o[12]
port 317 nsew signal output
rlabel metal2 s 51184 0 51240 400 6 wbs_dat_o[13]
port 318 nsew signal output
rlabel metal2 s 53872 0 53928 400 6 wbs_dat_o[14]
port 319 nsew signal output
rlabel metal2 s 56560 0 56616 400 6 wbs_dat_o[15]
port 320 nsew signal output
rlabel metal2 s 59248 0 59304 400 6 wbs_dat_o[16]
port 321 nsew signal output
rlabel metal2 s 61936 0 61992 400 6 wbs_dat_o[17]
port 322 nsew signal output
rlabel metal2 s 64624 0 64680 400 6 wbs_dat_o[18]
port 323 nsew signal output
rlabel metal2 s 67312 0 67368 400 6 wbs_dat_o[19]
port 324 nsew signal output
rlabel metal2 s 16240 0 16296 400 6 wbs_dat_o[1]
port 325 nsew signal output
rlabel metal2 s 70000 0 70056 400 6 wbs_dat_o[20]
port 326 nsew signal output
rlabel metal2 s 72688 0 72744 400 6 wbs_dat_o[21]
port 327 nsew signal output
rlabel metal2 s 75376 0 75432 400 6 wbs_dat_o[22]
port 328 nsew signal output
rlabel metal2 s 78064 0 78120 400 6 wbs_dat_o[23]
port 329 nsew signal output
rlabel metal2 s 80752 0 80808 400 6 wbs_dat_o[24]
port 330 nsew signal output
rlabel metal2 s 83440 0 83496 400 6 wbs_dat_o[25]
port 331 nsew signal output
rlabel metal2 s 86128 0 86184 400 6 wbs_dat_o[26]
port 332 nsew signal output
rlabel metal2 s 88816 0 88872 400 6 wbs_dat_o[27]
port 333 nsew signal output
rlabel metal2 s 91504 0 91560 400 6 wbs_dat_o[28]
port 334 nsew signal output
rlabel metal2 s 94192 0 94248 400 6 wbs_dat_o[29]
port 335 nsew signal output
rlabel metal2 s 19824 0 19880 400 6 wbs_dat_o[2]
port 336 nsew signal output
rlabel metal2 s 96880 0 96936 400 6 wbs_dat_o[30]
port 337 nsew signal output
rlabel metal2 s 99568 0 99624 400 6 wbs_dat_o[31]
port 338 nsew signal output
rlabel metal2 s 23408 0 23464 400 6 wbs_dat_o[3]
port 339 nsew signal output
rlabel metal2 s 26992 0 27048 400 6 wbs_dat_o[4]
port 340 nsew signal output
rlabel metal2 s 29680 0 29736 400 6 wbs_dat_o[5]
port 341 nsew signal output
rlabel metal2 s 32368 0 32424 400 6 wbs_dat_o[6]
port 342 nsew signal output
rlabel metal2 s 35056 0 35112 400 6 wbs_dat_o[7]
port 343 nsew signal output
rlabel metal2 s 37744 0 37800 400 6 wbs_dat_o[8]
port 344 nsew signal output
rlabel metal2 s 40432 0 40488 400 6 wbs_dat_o[9]
port 345 nsew signal output
rlabel metal2 s 13552 0 13608 400 6 wbs_sel_i[0]
port 346 nsew signal input
rlabel metal2 s 17136 0 17192 400 6 wbs_sel_i[1]
port 347 nsew signal input
rlabel metal2 s 20720 0 20776 400 6 wbs_sel_i[2]
port 348 nsew signal input
rlabel metal2 s 24304 0 24360 400 6 wbs_sel_i[3]
port 349 nsew signal input
rlabel metal2 s 9072 0 9128 400 6 wbs_stb_i
port 350 nsew signal input
rlabel metal2 s 9968 0 10024 400 6 wbs_we_i
port 351 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 280000 250000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 22296982
string GDS_FILE /home/navaneeth/Projects/openmpw/riscv_soc/openlane/user_proj_example/runs/23_11_30_17_09/results/signoff/user_proj_example.magic.gds
string GDS_START 284186
<< end >>


magic
tech gf180mcuD
magscale 1 5
timestamp 1701422585
<< obsm1 >>
rect 672 855 279328 174078
<< metal2 >>
rect 5936 175600 5992 176000
rect 16240 175600 16296 176000
rect 26544 175600 26600 176000
rect 36848 175600 36904 176000
rect 47152 175600 47208 176000
rect 57456 175600 57512 176000
rect 67760 175600 67816 176000
rect 78064 175600 78120 176000
rect 88368 175600 88424 176000
rect 98672 175600 98728 176000
rect 108976 175600 109032 176000
rect 119280 175600 119336 176000
rect 129584 175600 129640 176000
rect 139888 175600 139944 176000
rect 150192 175600 150248 176000
rect 160496 175600 160552 176000
rect 170800 175600 170856 176000
rect 181104 175600 181160 176000
rect 191408 175600 191464 176000
rect 201712 175600 201768 176000
rect 212016 175600 212072 176000
rect 222320 175600 222376 176000
rect 232624 175600 232680 176000
rect 242928 175600 242984 176000
rect 253232 175600 253288 176000
rect 263536 175600 263592 176000
rect 273840 175600 273896 176000
rect 5040 0 5096 400
rect 6608 0 6664 400
rect 8176 0 8232 400
rect 9744 0 9800 400
rect 11312 0 11368 400
rect 12880 0 12936 400
rect 14448 0 14504 400
rect 16016 0 16072 400
rect 17584 0 17640 400
rect 19152 0 19208 400
rect 20720 0 20776 400
rect 22288 0 22344 400
rect 23856 0 23912 400
rect 25424 0 25480 400
rect 26992 0 27048 400
rect 28560 0 28616 400
rect 30128 0 30184 400
rect 31696 0 31752 400
rect 33264 0 33320 400
rect 34832 0 34888 400
rect 36400 0 36456 400
rect 37968 0 38024 400
rect 39536 0 39592 400
rect 41104 0 41160 400
rect 42672 0 42728 400
rect 44240 0 44296 400
rect 45808 0 45864 400
rect 47376 0 47432 400
rect 48944 0 49000 400
rect 50512 0 50568 400
rect 52080 0 52136 400
rect 53648 0 53704 400
rect 55216 0 55272 400
rect 56784 0 56840 400
rect 58352 0 58408 400
rect 59920 0 59976 400
rect 61488 0 61544 400
rect 63056 0 63112 400
rect 64624 0 64680 400
rect 66192 0 66248 400
rect 67760 0 67816 400
rect 69328 0 69384 400
rect 70896 0 70952 400
rect 72464 0 72520 400
rect 74032 0 74088 400
rect 75600 0 75656 400
rect 77168 0 77224 400
rect 78736 0 78792 400
rect 80304 0 80360 400
rect 81872 0 81928 400
rect 83440 0 83496 400
rect 85008 0 85064 400
rect 86576 0 86632 400
rect 88144 0 88200 400
rect 89712 0 89768 400
rect 91280 0 91336 400
rect 92848 0 92904 400
rect 94416 0 94472 400
rect 95984 0 96040 400
rect 97552 0 97608 400
rect 99120 0 99176 400
rect 100688 0 100744 400
rect 102256 0 102312 400
rect 103824 0 103880 400
rect 105392 0 105448 400
rect 106960 0 107016 400
rect 108528 0 108584 400
rect 110096 0 110152 400
rect 111664 0 111720 400
rect 113232 0 113288 400
rect 114800 0 114856 400
rect 116368 0 116424 400
rect 117936 0 117992 400
rect 119504 0 119560 400
rect 121072 0 121128 400
rect 122640 0 122696 400
rect 124208 0 124264 400
rect 125776 0 125832 400
rect 127344 0 127400 400
rect 128912 0 128968 400
rect 130480 0 130536 400
rect 132048 0 132104 400
rect 133616 0 133672 400
rect 135184 0 135240 400
rect 136752 0 136808 400
rect 138320 0 138376 400
rect 139888 0 139944 400
rect 141456 0 141512 400
rect 143024 0 143080 400
rect 144592 0 144648 400
rect 146160 0 146216 400
rect 147728 0 147784 400
rect 149296 0 149352 400
rect 150864 0 150920 400
rect 152432 0 152488 400
rect 154000 0 154056 400
rect 155568 0 155624 400
rect 157136 0 157192 400
rect 158704 0 158760 400
rect 160272 0 160328 400
rect 161840 0 161896 400
rect 163408 0 163464 400
rect 164976 0 165032 400
rect 166544 0 166600 400
rect 168112 0 168168 400
rect 169680 0 169736 400
rect 171248 0 171304 400
rect 172816 0 172872 400
rect 174384 0 174440 400
rect 175952 0 176008 400
rect 177520 0 177576 400
rect 179088 0 179144 400
rect 180656 0 180712 400
rect 182224 0 182280 400
rect 183792 0 183848 400
rect 185360 0 185416 400
rect 186928 0 186984 400
rect 188496 0 188552 400
rect 190064 0 190120 400
rect 191632 0 191688 400
rect 193200 0 193256 400
rect 194768 0 194824 400
rect 196336 0 196392 400
rect 197904 0 197960 400
rect 199472 0 199528 400
rect 201040 0 201096 400
rect 202608 0 202664 400
rect 204176 0 204232 400
rect 205744 0 205800 400
rect 207312 0 207368 400
rect 208880 0 208936 400
rect 210448 0 210504 400
rect 212016 0 212072 400
rect 213584 0 213640 400
rect 215152 0 215208 400
rect 216720 0 216776 400
rect 218288 0 218344 400
rect 219856 0 219912 400
rect 221424 0 221480 400
rect 222992 0 223048 400
rect 224560 0 224616 400
rect 226128 0 226184 400
rect 227696 0 227752 400
rect 229264 0 229320 400
rect 230832 0 230888 400
rect 232400 0 232456 400
rect 233968 0 234024 400
rect 235536 0 235592 400
rect 237104 0 237160 400
rect 238672 0 238728 400
rect 240240 0 240296 400
rect 241808 0 241864 400
rect 243376 0 243432 400
rect 244944 0 245000 400
rect 246512 0 246568 400
rect 248080 0 248136 400
rect 249648 0 249704 400
rect 251216 0 251272 400
rect 252784 0 252840 400
rect 254352 0 254408 400
rect 255920 0 255976 400
rect 257488 0 257544 400
rect 259056 0 259112 400
rect 260624 0 260680 400
rect 262192 0 262248 400
rect 263760 0 263816 400
rect 265328 0 265384 400
rect 266896 0 266952 400
rect 268464 0 268520 400
rect 270032 0 270088 400
rect 271600 0 271656 400
rect 273168 0 273224 400
rect 274736 0 274792 400
<< obsm2 >>
rect 854 175570 5906 175658
rect 6022 175570 16210 175658
rect 16326 175570 26514 175658
rect 26630 175570 36818 175658
rect 36934 175570 47122 175658
rect 47238 175570 57426 175658
rect 57542 175570 67730 175658
rect 67846 175570 78034 175658
rect 78150 175570 88338 175658
rect 88454 175570 98642 175658
rect 98758 175570 108946 175658
rect 109062 175570 119250 175658
rect 119366 175570 129554 175658
rect 129670 175570 139858 175658
rect 139974 175570 150162 175658
rect 150278 175570 160466 175658
rect 160582 175570 170770 175658
rect 170886 175570 181074 175658
rect 181190 175570 191378 175658
rect 191494 175570 201682 175658
rect 201798 175570 211986 175658
rect 212102 175570 222290 175658
rect 222406 175570 232594 175658
rect 232710 175570 242898 175658
rect 243014 175570 253202 175658
rect 253318 175570 263506 175658
rect 263622 175570 273810 175658
rect 273926 175570 279146 175658
rect 854 430 279146 175570
rect 854 350 5010 430
rect 5126 350 6578 430
rect 6694 350 8146 430
rect 8262 350 9714 430
rect 9830 350 11282 430
rect 11398 350 12850 430
rect 12966 350 14418 430
rect 14534 350 15986 430
rect 16102 350 17554 430
rect 17670 350 19122 430
rect 19238 350 20690 430
rect 20806 350 22258 430
rect 22374 350 23826 430
rect 23942 350 25394 430
rect 25510 350 26962 430
rect 27078 350 28530 430
rect 28646 350 30098 430
rect 30214 350 31666 430
rect 31782 350 33234 430
rect 33350 350 34802 430
rect 34918 350 36370 430
rect 36486 350 37938 430
rect 38054 350 39506 430
rect 39622 350 41074 430
rect 41190 350 42642 430
rect 42758 350 44210 430
rect 44326 350 45778 430
rect 45894 350 47346 430
rect 47462 350 48914 430
rect 49030 350 50482 430
rect 50598 350 52050 430
rect 52166 350 53618 430
rect 53734 350 55186 430
rect 55302 350 56754 430
rect 56870 350 58322 430
rect 58438 350 59890 430
rect 60006 350 61458 430
rect 61574 350 63026 430
rect 63142 350 64594 430
rect 64710 350 66162 430
rect 66278 350 67730 430
rect 67846 350 69298 430
rect 69414 350 70866 430
rect 70982 350 72434 430
rect 72550 350 74002 430
rect 74118 350 75570 430
rect 75686 350 77138 430
rect 77254 350 78706 430
rect 78822 350 80274 430
rect 80390 350 81842 430
rect 81958 350 83410 430
rect 83526 350 84978 430
rect 85094 350 86546 430
rect 86662 350 88114 430
rect 88230 350 89682 430
rect 89798 350 91250 430
rect 91366 350 92818 430
rect 92934 350 94386 430
rect 94502 350 95954 430
rect 96070 350 97522 430
rect 97638 350 99090 430
rect 99206 350 100658 430
rect 100774 350 102226 430
rect 102342 350 103794 430
rect 103910 350 105362 430
rect 105478 350 106930 430
rect 107046 350 108498 430
rect 108614 350 110066 430
rect 110182 350 111634 430
rect 111750 350 113202 430
rect 113318 350 114770 430
rect 114886 350 116338 430
rect 116454 350 117906 430
rect 118022 350 119474 430
rect 119590 350 121042 430
rect 121158 350 122610 430
rect 122726 350 124178 430
rect 124294 350 125746 430
rect 125862 350 127314 430
rect 127430 350 128882 430
rect 128998 350 130450 430
rect 130566 350 132018 430
rect 132134 350 133586 430
rect 133702 350 135154 430
rect 135270 350 136722 430
rect 136838 350 138290 430
rect 138406 350 139858 430
rect 139974 350 141426 430
rect 141542 350 142994 430
rect 143110 350 144562 430
rect 144678 350 146130 430
rect 146246 350 147698 430
rect 147814 350 149266 430
rect 149382 350 150834 430
rect 150950 350 152402 430
rect 152518 350 153970 430
rect 154086 350 155538 430
rect 155654 350 157106 430
rect 157222 350 158674 430
rect 158790 350 160242 430
rect 160358 350 161810 430
rect 161926 350 163378 430
rect 163494 350 164946 430
rect 165062 350 166514 430
rect 166630 350 168082 430
rect 168198 350 169650 430
rect 169766 350 171218 430
rect 171334 350 172786 430
rect 172902 350 174354 430
rect 174470 350 175922 430
rect 176038 350 177490 430
rect 177606 350 179058 430
rect 179174 350 180626 430
rect 180742 350 182194 430
rect 182310 350 183762 430
rect 183878 350 185330 430
rect 185446 350 186898 430
rect 187014 350 188466 430
rect 188582 350 190034 430
rect 190150 350 191602 430
rect 191718 350 193170 430
rect 193286 350 194738 430
rect 194854 350 196306 430
rect 196422 350 197874 430
rect 197990 350 199442 430
rect 199558 350 201010 430
rect 201126 350 202578 430
rect 202694 350 204146 430
rect 204262 350 205714 430
rect 205830 350 207282 430
rect 207398 350 208850 430
rect 208966 350 210418 430
rect 210534 350 211986 430
rect 212102 350 213554 430
rect 213670 350 215122 430
rect 215238 350 216690 430
rect 216806 350 218258 430
rect 218374 350 219826 430
rect 219942 350 221394 430
rect 221510 350 222962 430
rect 223078 350 224530 430
rect 224646 350 226098 430
rect 226214 350 227666 430
rect 227782 350 229234 430
rect 229350 350 230802 430
rect 230918 350 232370 430
rect 232486 350 233938 430
rect 234054 350 235506 430
rect 235622 350 237074 430
rect 237190 350 238642 430
rect 238758 350 240210 430
rect 240326 350 241778 430
rect 241894 350 243346 430
rect 243462 350 244914 430
rect 245030 350 246482 430
rect 246598 350 248050 430
rect 248166 350 249618 430
rect 249734 350 251186 430
rect 251302 350 252754 430
rect 252870 350 254322 430
rect 254438 350 255890 430
rect 256006 350 257458 430
rect 257574 350 259026 430
rect 259142 350 260594 430
rect 260710 350 262162 430
rect 262278 350 263730 430
rect 263846 350 265298 430
rect 265414 350 266866 430
rect 266982 350 268434 430
rect 268550 350 270002 430
rect 270118 350 271570 430
rect 271686 350 273138 430
rect 273254 350 274706 430
rect 274822 350 279146 430
<< metal3 >>
rect 0 172928 400 172984
rect 279600 171696 280000 171752
rect 0 168784 400 168840
rect 279600 167888 280000 167944
rect 0 164640 400 164696
rect 279600 164080 280000 164136
rect 0 160496 400 160552
rect 279600 160272 280000 160328
rect 279600 156464 280000 156520
rect 0 156352 400 156408
rect 279600 152656 280000 152712
rect 0 152208 400 152264
rect 279600 148848 280000 148904
rect 0 148064 400 148120
rect 279600 145040 280000 145096
rect 0 143920 400 143976
rect 279600 141232 280000 141288
rect 0 139776 400 139832
rect 279600 137424 280000 137480
rect 0 135632 400 135688
rect 279600 133616 280000 133672
rect 0 131488 400 131544
rect 279600 129808 280000 129864
rect 0 127344 400 127400
rect 279600 126000 280000 126056
rect 0 123200 400 123256
rect 279600 122192 280000 122248
rect 0 119056 400 119112
rect 279600 118384 280000 118440
rect 0 114912 400 114968
rect 279600 114576 280000 114632
rect 0 110768 400 110824
rect 279600 110768 280000 110824
rect 279600 106960 280000 107016
rect 0 106624 400 106680
rect 279600 103152 280000 103208
rect 0 102480 400 102536
rect 279600 99344 280000 99400
rect 0 98336 400 98392
rect 279600 95536 280000 95592
rect 0 94192 400 94248
rect 279600 91728 280000 91784
rect 0 90048 400 90104
rect 279600 87920 280000 87976
rect 0 85904 400 85960
rect 279600 84112 280000 84168
rect 0 81760 400 81816
rect 279600 80304 280000 80360
rect 0 77616 400 77672
rect 279600 76496 280000 76552
rect 0 73472 400 73528
rect 279600 72688 280000 72744
rect 0 69328 400 69384
rect 279600 68880 280000 68936
rect 0 65184 400 65240
rect 279600 65072 280000 65128
rect 279600 61264 280000 61320
rect 0 61040 400 61096
rect 279600 57456 280000 57512
rect 0 56896 400 56952
rect 279600 53648 280000 53704
rect 0 52752 400 52808
rect 279600 49840 280000 49896
rect 0 48608 400 48664
rect 279600 46032 280000 46088
rect 0 44464 400 44520
rect 279600 42224 280000 42280
rect 0 40320 400 40376
rect 279600 38416 280000 38472
rect 0 36176 400 36232
rect 279600 34608 280000 34664
rect 0 32032 400 32088
rect 279600 30800 280000 30856
rect 0 27888 400 27944
rect 279600 26992 280000 27048
rect 0 23744 400 23800
rect 279600 23184 280000 23240
rect 0 19600 400 19656
rect 279600 19376 280000 19432
rect 279600 15568 280000 15624
rect 0 15456 400 15512
rect 279600 11760 280000 11816
rect 0 11312 400 11368
rect 279600 7952 280000 8008
rect 0 7168 400 7224
rect 279600 4144 280000 4200
rect 0 3024 400 3080
<< obsm3 >>
rect 400 173014 279650 174062
rect 430 172898 279650 173014
rect 400 171782 279650 172898
rect 400 171666 279570 171782
rect 400 168870 279650 171666
rect 430 168754 279650 168870
rect 400 167974 279650 168754
rect 400 167858 279570 167974
rect 400 164726 279650 167858
rect 430 164610 279650 164726
rect 400 164166 279650 164610
rect 400 164050 279570 164166
rect 400 160582 279650 164050
rect 430 160466 279650 160582
rect 400 160358 279650 160466
rect 400 160242 279570 160358
rect 400 156550 279650 160242
rect 400 156438 279570 156550
rect 430 156434 279570 156438
rect 430 156322 279650 156434
rect 400 152742 279650 156322
rect 400 152626 279570 152742
rect 400 152294 279650 152626
rect 430 152178 279650 152294
rect 400 148934 279650 152178
rect 400 148818 279570 148934
rect 400 148150 279650 148818
rect 430 148034 279650 148150
rect 400 145126 279650 148034
rect 400 145010 279570 145126
rect 400 144006 279650 145010
rect 430 143890 279650 144006
rect 400 141318 279650 143890
rect 400 141202 279570 141318
rect 400 139862 279650 141202
rect 430 139746 279650 139862
rect 400 137510 279650 139746
rect 400 137394 279570 137510
rect 400 135718 279650 137394
rect 430 135602 279650 135718
rect 400 133702 279650 135602
rect 400 133586 279570 133702
rect 400 131574 279650 133586
rect 430 131458 279650 131574
rect 400 129894 279650 131458
rect 400 129778 279570 129894
rect 400 127430 279650 129778
rect 430 127314 279650 127430
rect 400 126086 279650 127314
rect 400 125970 279570 126086
rect 400 123286 279650 125970
rect 430 123170 279650 123286
rect 400 122278 279650 123170
rect 400 122162 279570 122278
rect 400 119142 279650 122162
rect 430 119026 279650 119142
rect 400 118470 279650 119026
rect 400 118354 279570 118470
rect 400 114998 279650 118354
rect 430 114882 279650 114998
rect 400 114662 279650 114882
rect 400 114546 279570 114662
rect 400 110854 279650 114546
rect 430 110738 279570 110854
rect 400 107046 279650 110738
rect 400 106930 279570 107046
rect 400 106710 279650 106930
rect 430 106594 279650 106710
rect 400 103238 279650 106594
rect 400 103122 279570 103238
rect 400 102566 279650 103122
rect 430 102450 279650 102566
rect 400 99430 279650 102450
rect 400 99314 279570 99430
rect 400 98422 279650 99314
rect 430 98306 279650 98422
rect 400 95622 279650 98306
rect 400 95506 279570 95622
rect 400 94278 279650 95506
rect 430 94162 279650 94278
rect 400 91814 279650 94162
rect 400 91698 279570 91814
rect 400 90134 279650 91698
rect 430 90018 279650 90134
rect 400 88006 279650 90018
rect 400 87890 279570 88006
rect 400 85990 279650 87890
rect 430 85874 279650 85990
rect 400 84198 279650 85874
rect 400 84082 279570 84198
rect 400 81846 279650 84082
rect 430 81730 279650 81846
rect 400 80390 279650 81730
rect 400 80274 279570 80390
rect 400 77702 279650 80274
rect 430 77586 279650 77702
rect 400 76582 279650 77586
rect 400 76466 279570 76582
rect 400 73558 279650 76466
rect 430 73442 279650 73558
rect 400 72774 279650 73442
rect 400 72658 279570 72774
rect 400 69414 279650 72658
rect 430 69298 279650 69414
rect 400 68966 279650 69298
rect 400 68850 279570 68966
rect 400 65270 279650 68850
rect 430 65158 279650 65270
rect 430 65154 279570 65158
rect 400 65042 279570 65154
rect 400 61350 279650 65042
rect 400 61234 279570 61350
rect 400 61126 279650 61234
rect 430 61010 279650 61126
rect 400 57542 279650 61010
rect 400 57426 279570 57542
rect 400 56982 279650 57426
rect 430 56866 279650 56982
rect 400 53734 279650 56866
rect 400 53618 279570 53734
rect 400 52838 279650 53618
rect 430 52722 279650 52838
rect 400 49926 279650 52722
rect 400 49810 279570 49926
rect 400 48694 279650 49810
rect 430 48578 279650 48694
rect 400 46118 279650 48578
rect 400 46002 279570 46118
rect 400 44550 279650 46002
rect 430 44434 279650 44550
rect 400 42310 279650 44434
rect 400 42194 279570 42310
rect 400 40406 279650 42194
rect 430 40290 279650 40406
rect 400 38502 279650 40290
rect 400 38386 279570 38502
rect 400 36262 279650 38386
rect 430 36146 279650 36262
rect 400 34694 279650 36146
rect 400 34578 279570 34694
rect 400 32118 279650 34578
rect 430 32002 279650 32118
rect 400 30886 279650 32002
rect 400 30770 279570 30886
rect 400 27974 279650 30770
rect 430 27858 279650 27974
rect 400 27078 279650 27858
rect 400 26962 279570 27078
rect 400 23830 279650 26962
rect 430 23714 279650 23830
rect 400 23270 279650 23714
rect 400 23154 279570 23270
rect 400 19686 279650 23154
rect 430 19570 279650 19686
rect 400 19462 279650 19570
rect 400 19346 279570 19462
rect 400 15654 279650 19346
rect 400 15542 279570 15654
rect 430 15538 279570 15542
rect 430 15426 279650 15538
rect 400 11846 279650 15426
rect 400 11730 279570 11846
rect 400 11398 279650 11730
rect 430 11282 279650 11398
rect 400 8038 279650 11282
rect 400 7922 279570 8038
rect 400 7254 279650 7922
rect 430 7138 279650 7254
rect 400 4230 279650 7138
rect 400 4114 279570 4230
rect 400 3110 279650 4114
rect 430 2994 279650 3110
rect 400 1554 279650 2994
<< metal4 >>
rect 2224 1538 2384 174078
rect 9904 1538 10064 174078
rect 17584 1538 17744 174078
rect 25264 1538 25424 174078
rect 32944 1538 33104 174078
rect 40624 1538 40784 174078
rect 48304 1538 48464 174078
rect 55984 1538 56144 174078
rect 63664 1538 63824 174078
rect 71344 1538 71504 174078
rect 79024 1538 79184 174078
rect 86704 1538 86864 174078
rect 94384 1538 94544 174078
rect 102064 1538 102224 174078
rect 109744 1538 109904 174078
rect 117424 1538 117584 174078
rect 125104 1538 125264 174078
rect 132784 1538 132944 174078
rect 140464 1538 140624 174078
rect 148144 1538 148304 174078
rect 155824 1538 155984 174078
rect 163504 1538 163664 174078
rect 171184 1538 171344 174078
rect 178864 1538 179024 174078
rect 186544 1538 186704 174078
rect 194224 1538 194384 174078
rect 201904 1538 202064 174078
rect 209584 1538 209744 174078
rect 217264 1538 217424 174078
rect 224944 1538 225104 174078
rect 232624 1538 232784 174078
rect 240304 1538 240464 174078
rect 247984 1538 248144 174078
rect 255664 1538 255824 174078
rect 263344 1538 263504 174078
rect 271024 1538 271184 174078
rect 278704 1538 278864 174078
<< obsm4 >>
rect 11774 2865 17554 106055
rect 17774 2865 25234 106055
rect 25454 2865 32914 106055
rect 33134 2865 40594 106055
rect 40814 2865 48274 106055
rect 48494 2865 55954 106055
rect 56174 2865 63634 106055
rect 63854 2865 71314 106055
rect 71534 2865 78994 106055
rect 79214 2865 86674 106055
rect 86894 2865 94354 106055
rect 94574 2865 102034 106055
rect 102254 2865 109714 106055
rect 109934 2865 117394 106055
rect 117614 2865 125074 106055
rect 125294 2865 132754 106055
rect 132974 2865 140434 106055
rect 140654 2865 148114 106055
rect 148334 2865 155794 106055
rect 156014 2865 163474 106055
rect 163694 2865 171154 106055
rect 171374 2865 178834 106055
rect 179054 2865 186514 106055
rect 186734 2865 194194 106055
rect 194414 2865 201874 106055
rect 202094 2865 205282 106055
<< labels >>
rlabel metal3 s 279600 4144 280000 4200 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 279600 118384 280000 118440 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 279600 129808 280000 129864 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 279600 141232 280000 141288 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 279600 152656 280000 152712 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 279600 164080 280000 164136 6 io_in[14]
port 6 nsew signal input
rlabel metal2 s 273840 175600 273896 176000 6 io_in[15]
port 7 nsew signal input
rlabel metal2 s 242928 175600 242984 176000 6 io_in[16]
port 8 nsew signal input
rlabel metal2 s 212016 175600 212072 176000 6 io_in[17]
port 9 nsew signal input
rlabel metal2 s 181104 175600 181160 176000 6 io_in[18]
port 10 nsew signal input
rlabel metal2 s 150192 175600 150248 176000 6 io_in[19]
port 11 nsew signal input
rlabel metal3 s 279600 15568 280000 15624 6 io_in[1]
port 12 nsew signal input
rlabel metal2 s 119280 175600 119336 176000 6 io_in[20]
port 13 nsew signal input
rlabel metal2 s 88368 175600 88424 176000 6 io_in[21]
port 14 nsew signal input
rlabel metal2 s 57456 175600 57512 176000 6 io_in[22]
port 15 nsew signal input
rlabel metal2 s 26544 175600 26600 176000 6 io_in[23]
port 16 nsew signal input
rlabel metal3 s 0 172928 400 172984 6 io_in[24]
port 17 nsew signal input
rlabel metal3 s 0 160496 400 160552 6 io_in[25]
port 18 nsew signal input
rlabel metal3 s 0 148064 400 148120 6 io_in[26]
port 19 nsew signal input
rlabel metal3 s 0 135632 400 135688 6 io_in[27]
port 20 nsew signal input
rlabel metal3 s 0 123200 400 123256 6 io_in[28]
port 21 nsew signal input
rlabel metal3 s 0 110768 400 110824 6 io_in[29]
port 22 nsew signal input
rlabel metal3 s 279600 26992 280000 27048 6 io_in[2]
port 23 nsew signal input
rlabel metal3 s 0 98336 400 98392 6 io_in[30]
port 24 nsew signal input
rlabel metal3 s 0 85904 400 85960 6 io_in[31]
port 25 nsew signal input
rlabel metal3 s 0 73472 400 73528 6 io_in[32]
port 26 nsew signal input
rlabel metal3 s 0 61040 400 61096 6 io_in[33]
port 27 nsew signal input
rlabel metal3 s 0 48608 400 48664 6 io_in[34]
port 28 nsew signal input
rlabel metal3 s 0 36176 400 36232 6 io_in[35]
port 29 nsew signal input
rlabel metal3 s 0 23744 400 23800 6 io_in[36]
port 30 nsew signal input
rlabel metal3 s 0 11312 400 11368 6 io_in[37]
port 31 nsew signal input
rlabel metal3 s 279600 38416 280000 38472 6 io_in[3]
port 32 nsew signal input
rlabel metal3 s 279600 49840 280000 49896 6 io_in[4]
port 33 nsew signal input
rlabel metal3 s 279600 61264 280000 61320 6 io_in[5]
port 34 nsew signal input
rlabel metal3 s 279600 72688 280000 72744 6 io_in[6]
port 35 nsew signal input
rlabel metal3 s 279600 84112 280000 84168 6 io_in[7]
port 36 nsew signal input
rlabel metal3 s 279600 95536 280000 95592 6 io_in[8]
port 37 nsew signal input
rlabel metal3 s 279600 106960 280000 107016 6 io_in[9]
port 38 nsew signal input
rlabel metal3 s 279600 11760 280000 11816 6 io_oeb[0]
port 39 nsew signal output
rlabel metal3 s 279600 126000 280000 126056 6 io_oeb[10]
port 40 nsew signal output
rlabel metal3 s 279600 137424 280000 137480 6 io_oeb[11]
port 41 nsew signal output
rlabel metal3 s 279600 148848 280000 148904 6 io_oeb[12]
port 42 nsew signal output
rlabel metal3 s 279600 160272 280000 160328 6 io_oeb[13]
port 43 nsew signal output
rlabel metal3 s 279600 171696 280000 171752 6 io_oeb[14]
port 44 nsew signal output
rlabel metal2 s 253232 175600 253288 176000 6 io_oeb[15]
port 45 nsew signal output
rlabel metal2 s 222320 175600 222376 176000 6 io_oeb[16]
port 46 nsew signal output
rlabel metal2 s 191408 175600 191464 176000 6 io_oeb[17]
port 47 nsew signal output
rlabel metal2 s 160496 175600 160552 176000 6 io_oeb[18]
port 48 nsew signal output
rlabel metal2 s 129584 175600 129640 176000 6 io_oeb[19]
port 49 nsew signal output
rlabel metal3 s 279600 23184 280000 23240 6 io_oeb[1]
port 50 nsew signal output
rlabel metal2 s 98672 175600 98728 176000 6 io_oeb[20]
port 51 nsew signal output
rlabel metal2 s 67760 175600 67816 176000 6 io_oeb[21]
port 52 nsew signal output
rlabel metal2 s 36848 175600 36904 176000 6 io_oeb[22]
port 53 nsew signal output
rlabel metal2 s 5936 175600 5992 176000 6 io_oeb[23]
port 54 nsew signal output
rlabel metal3 s 0 164640 400 164696 6 io_oeb[24]
port 55 nsew signal output
rlabel metal3 s 0 152208 400 152264 6 io_oeb[25]
port 56 nsew signal output
rlabel metal3 s 0 139776 400 139832 6 io_oeb[26]
port 57 nsew signal output
rlabel metal3 s 0 127344 400 127400 6 io_oeb[27]
port 58 nsew signal output
rlabel metal3 s 0 114912 400 114968 6 io_oeb[28]
port 59 nsew signal output
rlabel metal3 s 0 102480 400 102536 6 io_oeb[29]
port 60 nsew signal output
rlabel metal3 s 279600 34608 280000 34664 6 io_oeb[2]
port 61 nsew signal output
rlabel metal3 s 0 90048 400 90104 6 io_oeb[30]
port 62 nsew signal output
rlabel metal3 s 0 77616 400 77672 6 io_oeb[31]
port 63 nsew signal output
rlabel metal3 s 0 65184 400 65240 6 io_oeb[32]
port 64 nsew signal output
rlabel metal3 s 0 52752 400 52808 6 io_oeb[33]
port 65 nsew signal output
rlabel metal3 s 0 40320 400 40376 6 io_oeb[34]
port 66 nsew signal output
rlabel metal3 s 0 27888 400 27944 6 io_oeb[35]
port 67 nsew signal output
rlabel metal3 s 0 15456 400 15512 6 io_oeb[36]
port 68 nsew signal output
rlabel metal3 s 0 3024 400 3080 6 io_oeb[37]
port 69 nsew signal output
rlabel metal3 s 279600 46032 280000 46088 6 io_oeb[3]
port 70 nsew signal output
rlabel metal3 s 279600 57456 280000 57512 6 io_oeb[4]
port 71 nsew signal output
rlabel metal3 s 279600 68880 280000 68936 6 io_oeb[5]
port 72 nsew signal output
rlabel metal3 s 279600 80304 280000 80360 6 io_oeb[6]
port 73 nsew signal output
rlabel metal3 s 279600 91728 280000 91784 6 io_oeb[7]
port 74 nsew signal output
rlabel metal3 s 279600 103152 280000 103208 6 io_oeb[8]
port 75 nsew signal output
rlabel metal3 s 279600 114576 280000 114632 6 io_oeb[9]
port 76 nsew signal output
rlabel metal3 s 279600 7952 280000 8008 6 io_out[0]
port 77 nsew signal output
rlabel metal3 s 279600 122192 280000 122248 6 io_out[10]
port 78 nsew signal output
rlabel metal3 s 279600 133616 280000 133672 6 io_out[11]
port 79 nsew signal output
rlabel metal3 s 279600 145040 280000 145096 6 io_out[12]
port 80 nsew signal output
rlabel metal3 s 279600 156464 280000 156520 6 io_out[13]
port 81 nsew signal output
rlabel metal3 s 279600 167888 280000 167944 6 io_out[14]
port 82 nsew signal output
rlabel metal2 s 263536 175600 263592 176000 6 io_out[15]
port 83 nsew signal output
rlabel metal2 s 232624 175600 232680 176000 6 io_out[16]
port 84 nsew signal output
rlabel metal2 s 201712 175600 201768 176000 6 io_out[17]
port 85 nsew signal output
rlabel metal2 s 170800 175600 170856 176000 6 io_out[18]
port 86 nsew signal output
rlabel metal2 s 139888 175600 139944 176000 6 io_out[19]
port 87 nsew signal output
rlabel metal3 s 279600 19376 280000 19432 6 io_out[1]
port 88 nsew signal output
rlabel metal2 s 108976 175600 109032 176000 6 io_out[20]
port 89 nsew signal output
rlabel metal2 s 78064 175600 78120 176000 6 io_out[21]
port 90 nsew signal output
rlabel metal2 s 47152 175600 47208 176000 6 io_out[22]
port 91 nsew signal output
rlabel metal2 s 16240 175600 16296 176000 6 io_out[23]
port 92 nsew signal output
rlabel metal3 s 0 168784 400 168840 6 io_out[24]
port 93 nsew signal output
rlabel metal3 s 0 156352 400 156408 6 io_out[25]
port 94 nsew signal output
rlabel metal3 s 0 143920 400 143976 6 io_out[26]
port 95 nsew signal output
rlabel metal3 s 0 131488 400 131544 6 io_out[27]
port 96 nsew signal output
rlabel metal3 s 0 119056 400 119112 6 io_out[28]
port 97 nsew signal output
rlabel metal3 s 0 106624 400 106680 6 io_out[29]
port 98 nsew signal output
rlabel metal3 s 279600 30800 280000 30856 6 io_out[2]
port 99 nsew signal output
rlabel metal3 s 0 94192 400 94248 6 io_out[30]
port 100 nsew signal output
rlabel metal3 s 0 81760 400 81816 6 io_out[31]
port 101 nsew signal output
rlabel metal3 s 0 69328 400 69384 6 io_out[32]
port 102 nsew signal output
rlabel metal3 s 0 56896 400 56952 6 io_out[33]
port 103 nsew signal output
rlabel metal3 s 0 44464 400 44520 6 io_out[34]
port 104 nsew signal output
rlabel metal3 s 0 32032 400 32088 6 io_out[35]
port 105 nsew signal output
rlabel metal3 s 0 19600 400 19656 6 io_out[36]
port 106 nsew signal output
rlabel metal3 s 0 7168 400 7224 6 io_out[37]
port 107 nsew signal output
rlabel metal3 s 279600 42224 280000 42280 6 io_out[3]
port 108 nsew signal output
rlabel metal3 s 279600 53648 280000 53704 6 io_out[4]
port 109 nsew signal output
rlabel metal3 s 279600 65072 280000 65128 6 io_out[5]
port 110 nsew signal output
rlabel metal3 s 279600 76496 280000 76552 6 io_out[6]
port 111 nsew signal output
rlabel metal3 s 279600 87920 280000 87976 6 io_out[7]
port 112 nsew signal output
rlabel metal3 s 279600 99344 280000 99400 6 io_out[8]
port 113 nsew signal output
rlabel metal3 s 279600 110768 280000 110824 6 io_out[9]
port 114 nsew signal output
rlabel metal2 s 171248 0 171304 400 6 la_data_out[0]
port 115 nsew signal output
rlabel metal2 s 186928 0 186984 400 6 la_data_out[10]
port 116 nsew signal output
rlabel metal2 s 188496 0 188552 400 6 la_data_out[11]
port 117 nsew signal output
rlabel metal2 s 190064 0 190120 400 6 la_data_out[12]
port 118 nsew signal output
rlabel metal2 s 191632 0 191688 400 6 la_data_out[13]
port 119 nsew signal output
rlabel metal2 s 193200 0 193256 400 6 la_data_out[14]
port 120 nsew signal output
rlabel metal2 s 194768 0 194824 400 6 la_data_out[15]
port 121 nsew signal output
rlabel metal2 s 196336 0 196392 400 6 la_data_out[16]
port 122 nsew signal output
rlabel metal2 s 197904 0 197960 400 6 la_data_out[17]
port 123 nsew signal output
rlabel metal2 s 199472 0 199528 400 6 la_data_out[18]
port 124 nsew signal output
rlabel metal2 s 201040 0 201096 400 6 la_data_out[19]
port 125 nsew signal output
rlabel metal2 s 172816 0 172872 400 6 la_data_out[1]
port 126 nsew signal output
rlabel metal2 s 202608 0 202664 400 6 la_data_out[20]
port 127 nsew signal output
rlabel metal2 s 204176 0 204232 400 6 la_data_out[21]
port 128 nsew signal output
rlabel metal2 s 205744 0 205800 400 6 la_data_out[22]
port 129 nsew signal output
rlabel metal2 s 207312 0 207368 400 6 la_data_out[23]
port 130 nsew signal output
rlabel metal2 s 208880 0 208936 400 6 la_data_out[24]
port 131 nsew signal output
rlabel metal2 s 210448 0 210504 400 6 la_data_out[25]
port 132 nsew signal output
rlabel metal2 s 212016 0 212072 400 6 la_data_out[26]
port 133 nsew signal output
rlabel metal2 s 213584 0 213640 400 6 la_data_out[27]
port 134 nsew signal output
rlabel metal2 s 215152 0 215208 400 6 la_data_out[28]
port 135 nsew signal output
rlabel metal2 s 216720 0 216776 400 6 la_data_out[29]
port 136 nsew signal output
rlabel metal2 s 174384 0 174440 400 6 la_data_out[2]
port 137 nsew signal output
rlabel metal2 s 218288 0 218344 400 6 la_data_out[30]
port 138 nsew signal output
rlabel metal2 s 219856 0 219912 400 6 la_data_out[31]
port 139 nsew signal output
rlabel metal2 s 221424 0 221480 400 6 la_data_out[32]
port 140 nsew signal output
rlabel metal2 s 222992 0 223048 400 6 la_data_out[33]
port 141 nsew signal output
rlabel metal2 s 224560 0 224616 400 6 la_data_out[34]
port 142 nsew signal output
rlabel metal2 s 226128 0 226184 400 6 la_data_out[35]
port 143 nsew signal output
rlabel metal2 s 227696 0 227752 400 6 la_data_out[36]
port 144 nsew signal output
rlabel metal2 s 229264 0 229320 400 6 la_data_out[37]
port 145 nsew signal output
rlabel metal2 s 230832 0 230888 400 6 la_data_out[38]
port 146 nsew signal output
rlabel metal2 s 232400 0 232456 400 6 la_data_out[39]
port 147 nsew signal output
rlabel metal2 s 175952 0 176008 400 6 la_data_out[3]
port 148 nsew signal output
rlabel metal2 s 233968 0 234024 400 6 la_data_out[40]
port 149 nsew signal output
rlabel metal2 s 235536 0 235592 400 6 la_data_out[41]
port 150 nsew signal output
rlabel metal2 s 237104 0 237160 400 6 la_data_out[42]
port 151 nsew signal output
rlabel metal2 s 238672 0 238728 400 6 la_data_out[43]
port 152 nsew signal output
rlabel metal2 s 240240 0 240296 400 6 la_data_out[44]
port 153 nsew signal output
rlabel metal2 s 241808 0 241864 400 6 la_data_out[45]
port 154 nsew signal output
rlabel metal2 s 243376 0 243432 400 6 la_data_out[46]
port 155 nsew signal output
rlabel metal2 s 244944 0 245000 400 6 la_data_out[47]
port 156 nsew signal output
rlabel metal2 s 246512 0 246568 400 6 la_data_out[48]
port 157 nsew signal output
rlabel metal2 s 248080 0 248136 400 6 la_data_out[49]
port 158 nsew signal output
rlabel metal2 s 177520 0 177576 400 6 la_data_out[4]
port 159 nsew signal output
rlabel metal2 s 249648 0 249704 400 6 la_data_out[50]
port 160 nsew signal output
rlabel metal2 s 251216 0 251272 400 6 la_data_out[51]
port 161 nsew signal output
rlabel metal2 s 252784 0 252840 400 6 la_data_out[52]
port 162 nsew signal output
rlabel metal2 s 254352 0 254408 400 6 la_data_out[53]
port 163 nsew signal output
rlabel metal2 s 255920 0 255976 400 6 la_data_out[54]
port 164 nsew signal output
rlabel metal2 s 257488 0 257544 400 6 la_data_out[55]
port 165 nsew signal output
rlabel metal2 s 259056 0 259112 400 6 la_data_out[56]
port 166 nsew signal output
rlabel metal2 s 260624 0 260680 400 6 la_data_out[57]
port 167 nsew signal output
rlabel metal2 s 262192 0 262248 400 6 la_data_out[58]
port 168 nsew signal output
rlabel metal2 s 263760 0 263816 400 6 la_data_out[59]
port 169 nsew signal output
rlabel metal2 s 179088 0 179144 400 6 la_data_out[5]
port 170 nsew signal output
rlabel metal2 s 265328 0 265384 400 6 la_data_out[60]
port 171 nsew signal output
rlabel metal2 s 266896 0 266952 400 6 la_data_out[61]
port 172 nsew signal output
rlabel metal2 s 268464 0 268520 400 6 la_data_out[62]
port 173 nsew signal output
rlabel metal2 s 270032 0 270088 400 6 la_data_out[63]
port 174 nsew signal output
rlabel metal2 s 180656 0 180712 400 6 la_data_out[6]
port 175 nsew signal output
rlabel metal2 s 182224 0 182280 400 6 la_data_out[7]
port 176 nsew signal output
rlabel metal2 s 183792 0 183848 400 6 la_data_out[8]
port 177 nsew signal output
rlabel metal2 s 185360 0 185416 400 6 la_data_out[9]
port 178 nsew signal output
rlabel metal2 s 271600 0 271656 400 6 user_irq[0]
port 179 nsew signal output
rlabel metal2 s 273168 0 273224 400 6 user_irq[1]
port 180 nsew signal output
rlabel metal2 s 274736 0 274792 400 6 user_irq[2]
port 181 nsew signal output
rlabel metal4 s 2224 1538 2384 174078 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 174078 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 174078 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 174078 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 174078 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 174078 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 174078 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 109744 1538 109904 174078 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 125104 1538 125264 174078 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 140464 1538 140624 174078 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 155824 1538 155984 174078 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 171184 1538 171344 174078 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 186544 1538 186704 174078 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 201904 1538 202064 174078 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 217264 1538 217424 174078 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 232624 1538 232784 174078 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 247984 1538 248144 174078 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 263344 1538 263504 174078 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 278704 1538 278864 174078 6 vdd
port 182 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 174078 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 174078 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 174078 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 174078 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 174078 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 174078 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 174078 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 117424 1538 117584 174078 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 132784 1538 132944 174078 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 148144 1538 148304 174078 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 163504 1538 163664 174078 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 178864 1538 179024 174078 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 194224 1538 194384 174078 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 209584 1538 209744 174078 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 224944 1538 225104 174078 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 240304 1538 240464 174078 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 255664 1538 255824 174078 6 vss
port 183 nsew ground bidirectional
rlabel metal4 s 271024 1538 271184 174078 6 vss
port 183 nsew ground bidirectional
rlabel metal2 s 5040 0 5096 400 6 wb_clk_i
port 184 nsew signal input
rlabel metal2 s 6608 0 6664 400 6 wb_rst_i
port 185 nsew signal input
rlabel metal2 s 8176 0 8232 400 6 wbs_ack_o
port 186 nsew signal output
rlabel metal2 s 14448 0 14504 400 6 wbs_adr_i[0]
port 187 nsew signal input
rlabel metal2 s 67760 0 67816 400 6 wbs_adr_i[10]
port 188 nsew signal input
rlabel metal2 s 72464 0 72520 400 6 wbs_adr_i[11]
port 189 nsew signal input
rlabel metal2 s 77168 0 77224 400 6 wbs_adr_i[12]
port 190 nsew signal input
rlabel metal2 s 81872 0 81928 400 6 wbs_adr_i[13]
port 191 nsew signal input
rlabel metal2 s 86576 0 86632 400 6 wbs_adr_i[14]
port 192 nsew signal input
rlabel metal2 s 91280 0 91336 400 6 wbs_adr_i[15]
port 193 nsew signal input
rlabel metal2 s 95984 0 96040 400 6 wbs_adr_i[16]
port 194 nsew signal input
rlabel metal2 s 100688 0 100744 400 6 wbs_adr_i[17]
port 195 nsew signal input
rlabel metal2 s 105392 0 105448 400 6 wbs_adr_i[18]
port 196 nsew signal input
rlabel metal2 s 110096 0 110152 400 6 wbs_adr_i[19]
port 197 nsew signal input
rlabel metal2 s 20720 0 20776 400 6 wbs_adr_i[1]
port 198 nsew signal input
rlabel metal2 s 114800 0 114856 400 6 wbs_adr_i[20]
port 199 nsew signal input
rlabel metal2 s 119504 0 119560 400 6 wbs_adr_i[21]
port 200 nsew signal input
rlabel metal2 s 124208 0 124264 400 6 wbs_adr_i[22]
port 201 nsew signal input
rlabel metal2 s 128912 0 128968 400 6 wbs_adr_i[23]
port 202 nsew signal input
rlabel metal2 s 133616 0 133672 400 6 wbs_adr_i[24]
port 203 nsew signal input
rlabel metal2 s 138320 0 138376 400 6 wbs_adr_i[25]
port 204 nsew signal input
rlabel metal2 s 143024 0 143080 400 6 wbs_adr_i[26]
port 205 nsew signal input
rlabel metal2 s 147728 0 147784 400 6 wbs_adr_i[27]
port 206 nsew signal input
rlabel metal2 s 152432 0 152488 400 6 wbs_adr_i[28]
port 207 nsew signal input
rlabel metal2 s 157136 0 157192 400 6 wbs_adr_i[29]
port 208 nsew signal input
rlabel metal2 s 26992 0 27048 400 6 wbs_adr_i[2]
port 209 nsew signal input
rlabel metal2 s 161840 0 161896 400 6 wbs_adr_i[30]
port 210 nsew signal input
rlabel metal2 s 166544 0 166600 400 6 wbs_adr_i[31]
port 211 nsew signal input
rlabel metal2 s 33264 0 33320 400 6 wbs_adr_i[3]
port 212 nsew signal input
rlabel metal2 s 39536 0 39592 400 6 wbs_adr_i[4]
port 213 nsew signal input
rlabel metal2 s 44240 0 44296 400 6 wbs_adr_i[5]
port 214 nsew signal input
rlabel metal2 s 48944 0 49000 400 6 wbs_adr_i[6]
port 215 nsew signal input
rlabel metal2 s 53648 0 53704 400 6 wbs_adr_i[7]
port 216 nsew signal input
rlabel metal2 s 58352 0 58408 400 6 wbs_adr_i[8]
port 217 nsew signal input
rlabel metal2 s 63056 0 63112 400 6 wbs_adr_i[9]
port 218 nsew signal input
rlabel metal2 s 9744 0 9800 400 6 wbs_cyc_i
port 219 nsew signal input
rlabel metal2 s 16016 0 16072 400 6 wbs_dat_i[0]
port 220 nsew signal input
rlabel metal2 s 69328 0 69384 400 6 wbs_dat_i[10]
port 221 nsew signal input
rlabel metal2 s 74032 0 74088 400 6 wbs_dat_i[11]
port 222 nsew signal input
rlabel metal2 s 78736 0 78792 400 6 wbs_dat_i[12]
port 223 nsew signal input
rlabel metal2 s 83440 0 83496 400 6 wbs_dat_i[13]
port 224 nsew signal input
rlabel metal2 s 88144 0 88200 400 6 wbs_dat_i[14]
port 225 nsew signal input
rlabel metal2 s 92848 0 92904 400 6 wbs_dat_i[15]
port 226 nsew signal input
rlabel metal2 s 97552 0 97608 400 6 wbs_dat_i[16]
port 227 nsew signal input
rlabel metal2 s 102256 0 102312 400 6 wbs_dat_i[17]
port 228 nsew signal input
rlabel metal2 s 106960 0 107016 400 6 wbs_dat_i[18]
port 229 nsew signal input
rlabel metal2 s 111664 0 111720 400 6 wbs_dat_i[19]
port 230 nsew signal input
rlabel metal2 s 22288 0 22344 400 6 wbs_dat_i[1]
port 231 nsew signal input
rlabel metal2 s 116368 0 116424 400 6 wbs_dat_i[20]
port 232 nsew signal input
rlabel metal2 s 121072 0 121128 400 6 wbs_dat_i[21]
port 233 nsew signal input
rlabel metal2 s 125776 0 125832 400 6 wbs_dat_i[22]
port 234 nsew signal input
rlabel metal2 s 130480 0 130536 400 6 wbs_dat_i[23]
port 235 nsew signal input
rlabel metal2 s 135184 0 135240 400 6 wbs_dat_i[24]
port 236 nsew signal input
rlabel metal2 s 139888 0 139944 400 6 wbs_dat_i[25]
port 237 nsew signal input
rlabel metal2 s 144592 0 144648 400 6 wbs_dat_i[26]
port 238 nsew signal input
rlabel metal2 s 149296 0 149352 400 6 wbs_dat_i[27]
port 239 nsew signal input
rlabel metal2 s 154000 0 154056 400 6 wbs_dat_i[28]
port 240 nsew signal input
rlabel metal2 s 158704 0 158760 400 6 wbs_dat_i[29]
port 241 nsew signal input
rlabel metal2 s 28560 0 28616 400 6 wbs_dat_i[2]
port 242 nsew signal input
rlabel metal2 s 163408 0 163464 400 6 wbs_dat_i[30]
port 243 nsew signal input
rlabel metal2 s 168112 0 168168 400 6 wbs_dat_i[31]
port 244 nsew signal input
rlabel metal2 s 34832 0 34888 400 6 wbs_dat_i[3]
port 245 nsew signal input
rlabel metal2 s 41104 0 41160 400 6 wbs_dat_i[4]
port 246 nsew signal input
rlabel metal2 s 45808 0 45864 400 6 wbs_dat_i[5]
port 247 nsew signal input
rlabel metal2 s 50512 0 50568 400 6 wbs_dat_i[6]
port 248 nsew signal input
rlabel metal2 s 55216 0 55272 400 6 wbs_dat_i[7]
port 249 nsew signal input
rlabel metal2 s 59920 0 59976 400 6 wbs_dat_i[8]
port 250 nsew signal input
rlabel metal2 s 64624 0 64680 400 6 wbs_dat_i[9]
port 251 nsew signal input
rlabel metal2 s 17584 0 17640 400 6 wbs_dat_o[0]
port 252 nsew signal output
rlabel metal2 s 70896 0 70952 400 6 wbs_dat_o[10]
port 253 nsew signal output
rlabel metal2 s 75600 0 75656 400 6 wbs_dat_o[11]
port 254 nsew signal output
rlabel metal2 s 80304 0 80360 400 6 wbs_dat_o[12]
port 255 nsew signal output
rlabel metal2 s 85008 0 85064 400 6 wbs_dat_o[13]
port 256 nsew signal output
rlabel metal2 s 89712 0 89768 400 6 wbs_dat_o[14]
port 257 nsew signal output
rlabel metal2 s 94416 0 94472 400 6 wbs_dat_o[15]
port 258 nsew signal output
rlabel metal2 s 99120 0 99176 400 6 wbs_dat_o[16]
port 259 nsew signal output
rlabel metal2 s 103824 0 103880 400 6 wbs_dat_o[17]
port 260 nsew signal output
rlabel metal2 s 108528 0 108584 400 6 wbs_dat_o[18]
port 261 nsew signal output
rlabel metal2 s 113232 0 113288 400 6 wbs_dat_o[19]
port 262 nsew signal output
rlabel metal2 s 23856 0 23912 400 6 wbs_dat_o[1]
port 263 nsew signal output
rlabel metal2 s 117936 0 117992 400 6 wbs_dat_o[20]
port 264 nsew signal output
rlabel metal2 s 122640 0 122696 400 6 wbs_dat_o[21]
port 265 nsew signal output
rlabel metal2 s 127344 0 127400 400 6 wbs_dat_o[22]
port 266 nsew signal output
rlabel metal2 s 132048 0 132104 400 6 wbs_dat_o[23]
port 267 nsew signal output
rlabel metal2 s 136752 0 136808 400 6 wbs_dat_o[24]
port 268 nsew signal output
rlabel metal2 s 141456 0 141512 400 6 wbs_dat_o[25]
port 269 nsew signal output
rlabel metal2 s 146160 0 146216 400 6 wbs_dat_o[26]
port 270 nsew signal output
rlabel metal2 s 150864 0 150920 400 6 wbs_dat_o[27]
port 271 nsew signal output
rlabel metal2 s 155568 0 155624 400 6 wbs_dat_o[28]
port 272 nsew signal output
rlabel metal2 s 160272 0 160328 400 6 wbs_dat_o[29]
port 273 nsew signal output
rlabel metal2 s 30128 0 30184 400 6 wbs_dat_o[2]
port 274 nsew signal output
rlabel metal2 s 164976 0 165032 400 6 wbs_dat_o[30]
port 275 nsew signal output
rlabel metal2 s 169680 0 169736 400 6 wbs_dat_o[31]
port 276 nsew signal output
rlabel metal2 s 36400 0 36456 400 6 wbs_dat_o[3]
port 277 nsew signal output
rlabel metal2 s 42672 0 42728 400 6 wbs_dat_o[4]
port 278 nsew signal output
rlabel metal2 s 47376 0 47432 400 6 wbs_dat_o[5]
port 279 nsew signal output
rlabel metal2 s 52080 0 52136 400 6 wbs_dat_o[6]
port 280 nsew signal output
rlabel metal2 s 56784 0 56840 400 6 wbs_dat_o[7]
port 281 nsew signal output
rlabel metal2 s 61488 0 61544 400 6 wbs_dat_o[8]
port 282 nsew signal output
rlabel metal2 s 66192 0 66248 400 6 wbs_dat_o[9]
port 283 nsew signal output
rlabel metal2 s 19152 0 19208 400 6 wbs_sel_i[0]
port 284 nsew signal input
rlabel metal2 s 25424 0 25480 400 6 wbs_sel_i[1]
port 285 nsew signal input
rlabel metal2 s 31696 0 31752 400 6 wbs_sel_i[2]
port 286 nsew signal input
rlabel metal2 s 37968 0 38024 400 6 wbs_sel_i[3]
port 287 nsew signal input
rlabel metal2 s 11312 0 11368 400 6 wbs_stb_i
port 288 nsew signal input
rlabel metal2 s 12880 0 12936 400 6 wbs_we_i
port 289 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 280000 176000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 52216222
string GDS_FILE /home/navaneeth/Projects/openmpw/riscv_soc/openlane/alpha_soc/runs/23_12_01_14_26/results/signoff/alpha_soc.magic.gds
string GDS_START 554862
<< end >>

